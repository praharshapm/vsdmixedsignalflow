magic
tech sky130A
magscale 1 2
timestamp 1598265745
<< locali >>
rect 12541 2907 12575 3009
<< viali >>
rect 23765 27421 23799 27455
rect 23121 27353 23155 27387
rect 23213 27081 23247 27115
rect 16773 16677 16807 16711
rect 14197 16541 14231 16575
rect 16129 16541 16163 16575
rect 16497 16541 16531 16575
rect 16865 16541 16899 16575
rect 14381 16405 14415 16439
rect 15577 16405 15611 16439
rect 14197 16201 14231 16235
rect 16773 16201 16807 16235
rect 14749 16133 14783 16167
rect 14473 16065 14507 16099
rect 19901 16065 19935 16099
rect 16497 15997 16531 16031
rect 19257 15997 19291 16031
rect 13829 15861 13863 15895
rect 17141 15861 17175 15895
rect 16497 15657 16531 15691
rect 17417 15657 17451 15691
rect 14381 15521 14415 15555
rect 18061 15521 18095 15555
rect 19717 15521 19751 15555
rect 20085 15521 20119 15555
rect 23121 15521 23155 15555
rect 12817 15453 12851 15487
rect 14013 15453 14047 15487
rect 16129 15453 16163 15487
rect 17601 15453 17635 15487
rect 17785 15453 17819 15487
rect 18153 15453 18187 15487
rect 19165 15453 19199 15487
rect 21097 15453 21131 15487
rect 13553 15385 13587 15419
rect 13829 15385 13863 15419
rect 21373 15385 21407 15419
rect 13001 15317 13035 15351
rect 14657 15317 14691 15351
rect 15945 15317 15979 15351
rect 19349 15317 19383 15351
rect 12081 15113 12115 15147
rect 14933 15113 14967 15147
rect 21005 15113 21039 15147
rect 21649 15113 21683 15147
rect 21925 15113 21959 15147
rect 17601 15045 17635 15079
rect 18521 15045 18555 15079
rect 14657 14977 14691 15011
rect 15485 14977 15519 15011
rect 19441 14977 19475 15011
rect 19993 14977 20027 15011
rect 20177 14977 20211 15011
rect 21465 14977 21499 15011
rect 12633 14909 12667 14943
rect 12909 14909 12943 14943
rect 16497 14909 16531 14943
rect 19257 14909 19291 14943
rect 20545 14909 20579 14943
rect 16865 14841 16899 14875
rect 15669 14773 15703 14807
rect 17233 14773 17267 14807
rect 18889 14773 18923 14807
rect 14657 14569 14691 14603
rect 17417 14569 17451 14603
rect 18429 14569 18463 14603
rect 20269 14569 20303 14603
rect 21189 14569 21223 14603
rect 21557 14569 21591 14603
rect 12265 14433 12299 14467
rect 12909 14433 12943 14467
rect 14197 14433 14231 14467
rect 15577 14433 15611 14467
rect 16497 14433 16531 14467
rect 19257 14433 19291 14467
rect 22385 14433 22419 14467
rect 24409 14433 24443 14467
rect 11897 14365 11931 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 13737 14365 13771 14399
rect 14289 14365 14323 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 17601 14365 17635 14399
rect 18153 14365 18187 14399
rect 19441 14365 19475 14399
rect 19809 14365 19843 14399
rect 19993 14365 20027 14399
rect 16221 14297 16255 14331
rect 22661 14297 22695 14331
rect 12541 14229 12575 14263
rect 19073 14229 19107 14263
rect 12725 14025 12759 14059
rect 13093 14025 13127 14059
rect 15117 14025 15151 14059
rect 18981 14025 19015 14059
rect 20177 14025 20211 14059
rect 21465 14025 21499 14059
rect 23121 14025 23155 14059
rect 12081 13957 12115 13991
rect 13553 13957 13587 13991
rect 15577 13957 15611 13991
rect 17049 13957 17083 13991
rect 17693 13957 17727 13991
rect 8769 13889 8803 13923
rect 14013 13889 14047 13923
rect 14381 13889 14415 13923
rect 14473 13889 14507 13923
rect 15669 13889 15703 13923
rect 19349 13889 19383 13923
rect 19717 13889 19751 13923
rect 21005 13889 21039 13923
rect 21281 13889 21315 13923
rect 15393 13821 15427 13855
rect 16497 13821 16531 13855
rect 19165 13821 19199 13855
rect 19257 13821 19291 13855
rect 19625 13821 19659 13855
rect 20545 13821 20579 13855
rect 21097 13821 21131 13855
rect 22385 13753 22419 13787
rect 8953 13685 8987 13719
rect 11345 13685 11379 13719
rect 11713 13685 11747 13719
rect 15853 13685 15887 13719
rect 18429 13685 18463 13719
rect 22753 13685 22787 13719
rect 11529 13481 11563 13515
rect 12265 13481 12299 13515
rect 15761 13481 15795 13515
rect 18245 13481 18279 13515
rect 20085 13481 20119 13515
rect 20545 13481 20579 13515
rect 21557 13481 21591 13515
rect 12633 13413 12667 13447
rect 14749 13413 14783 13447
rect 18981 13413 19015 13447
rect 19625 13413 19659 13447
rect 21281 13413 21315 13447
rect 13001 13345 13035 13379
rect 13461 13345 13495 13379
rect 14197 13345 14231 13379
rect 15853 13345 15887 13379
rect 17049 13345 17083 13379
rect 13829 13277 13863 13311
rect 14105 13277 14139 13311
rect 15632 13277 15666 13311
rect 17141 13277 17175 13311
rect 19165 13277 19199 13311
rect 21097 13277 21131 13311
rect 15485 13209 15519 13243
rect 16773 13209 16807 13243
rect 17601 13209 17635 13243
rect 8769 13141 8803 13175
rect 11897 13141 11931 13175
rect 16129 13141 16163 13175
rect 23765 13141 23799 13175
rect 11621 12937 11655 12971
rect 15485 12937 15519 12971
rect 18521 12937 18555 12971
rect 19073 12937 19107 12971
rect 19533 12937 19567 12971
rect 18245 12869 18279 12903
rect 9137 12801 9171 12835
rect 13093 12801 13127 12835
rect 13277 12801 13311 12835
rect 13461 12801 13495 12835
rect 14013 12801 14047 12835
rect 16589 12801 16623 12835
rect 16865 12801 16899 12835
rect 18429 12801 18463 12835
rect 19901 12801 19935 12835
rect 20729 12801 20763 12835
rect 22017 12801 22051 12835
rect 22293 12801 22327 12835
rect 8677 12733 8711 12767
rect 12633 12733 12667 12767
rect 13737 12733 13771 12767
rect 16129 12733 16163 12767
rect 20453 12733 20487 12767
rect 20913 12733 20947 12767
rect 22385 12733 22419 12767
rect 16865 12665 16899 12699
rect 25329 12665 25363 12699
rect 12081 12597 12115 12631
rect 14381 12597 14415 12631
rect 14841 12597 14875 12631
rect 17509 12597 17543 12631
rect 21189 12597 21223 12631
rect 23213 12597 23247 12631
rect 9137 12393 9171 12427
rect 11253 12393 11287 12427
rect 13829 12393 13863 12427
rect 14289 12393 14323 12427
rect 17049 12393 17083 12427
rect 17693 12393 17727 12427
rect 19073 12393 19107 12427
rect 20269 12393 20303 12427
rect 24409 12393 24443 12427
rect 15945 12325 15979 12359
rect 18337 12325 18371 12359
rect 21281 12325 21315 12359
rect 22201 12325 22235 12359
rect 25145 12325 25179 12359
rect 8217 12257 8251 12291
rect 11805 12257 11839 12291
rect 15485 12257 15519 12291
rect 17417 12257 17451 12291
rect 8309 12189 8343 12223
rect 11529 12189 11563 12223
rect 16221 12189 16255 12223
rect 16497 12189 16531 12223
rect 17509 12189 17543 12223
rect 18981 12189 19015 12223
rect 21097 12189 21131 12223
rect 22385 12189 22419 12223
rect 22569 12189 22603 12223
rect 22753 12189 22787 12223
rect 8769 12121 8803 12155
rect 13553 12121 13587 12155
rect 18797 12121 18831 12155
rect 23213 12121 23247 12155
rect 10885 12053 10919 12087
rect 14933 12053 14967 12087
rect 19993 12053 20027 12087
rect 21649 12053 21683 12087
rect 8217 11849 8251 11883
rect 8585 11849 8619 11883
rect 10701 11849 10735 11883
rect 11529 11849 11563 11883
rect 13185 11849 13219 11883
rect 13645 11849 13679 11883
rect 14105 11849 14139 11883
rect 16589 11849 16623 11883
rect 17141 11849 17175 11883
rect 17417 11849 17451 11883
rect 18245 11849 18279 11883
rect 20453 11849 20487 11883
rect 22753 11849 22787 11883
rect 11069 11781 11103 11815
rect 21005 11781 21039 11815
rect 23121 11781 23155 11815
rect 9781 11713 9815 11747
rect 11345 11713 11379 11747
rect 12633 11713 12667 11747
rect 14933 11713 14967 11747
rect 15117 11713 15151 11747
rect 15209 11713 15243 11747
rect 15853 11713 15887 11747
rect 16957 11713 16991 11747
rect 18981 11713 19015 11747
rect 19441 11713 19475 11747
rect 19533 11713 19567 11747
rect 21741 11713 21775 11747
rect 22385 11713 22419 11747
rect 8953 11645 8987 11679
rect 9505 11645 9539 11679
rect 9965 11645 9999 11679
rect 14381 11645 14415 11679
rect 15669 11645 15703 11679
rect 18797 11645 18831 11679
rect 21373 11645 21407 11679
rect 12817 11577 12851 11611
rect 21281 11577 21315 11611
rect 11805 11509 11839 11543
rect 16221 11509 16255 11543
rect 19993 11509 20027 11543
rect 21143 11509 21177 11543
rect 22017 11509 22051 11543
rect 8677 11305 8711 11339
rect 12909 11305 12943 11339
rect 13277 11305 13311 11339
rect 13737 11305 13771 11339
rect 15577 11305 15611 11339
rect 19717 11305 19751 11339
rect 20453 11305 20487 11339
rect 22017 11305 22051 11339
rect 22937 11305 22971 11339
rect 9045 11237 9079 11271
rect 14841 11237 14875 11271
rect 22569 11237 22603 11271
rect 12081 11169 12115 11203
rect 16037 11169 16071 11203
rect 16589 11169 16623 11203
rect 18245 11169 18279 11203
rect 11253 11101 11287 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 12173 11101 12207 11135
rect 16129 11101 16163 11135
rect 16497 11101 16531 11135
rect 17785 11101 17819 11135
rect 18153 11101 18187 11135
rect 19349 11101 19383 11135
rect 21649 11101 21683 11135
rect 10793 11033 10827 11067
rect 14105 11033 14139 11067
rect 17325 11033 17359 11067
rect 8309 10965 8343 10999
rect 10425 10965 10459 10999
rect 12541 10965 12575 10999
rect 14381 10965 14415 10999
rect 17049 10965 17083 10999
rect 18797 10965 18831 10999
rect 21097 10965 21131 10999
rect 9781 10761 9815 10795
rect 11253 10761 11287 10795
rect 12725 10761 12759 10795
rect 13093 10761 13127 10795
rect 13461 10761 13495 10795
rect 16037 10761 16071 10795
rect 17509 10761 17543 10795
rect 19349 10761 19383 10795
rect 19625 10761 19659 10795
rect 22017 10761 22051 10795
rect 22385 10761 22419 10795
rect 22753 10761 22787 10795
rect 10885 10693 10919 10727
rect 15761 10693 15795 10727
rect 18981 10693 19015 10727
rect 20177 10693 20211 10727
rect 7665 10625 7699 10659
rect 8309 10625 8343 10659
rect 8769 10625 8803 10659
rect 9229 10625 9263 10659
rect 9321 10625 9355 10659
rect 11529 10625 11563 10659
rect 16957 10625 16991 10659
rect 18889 10625 18923 10659
rect 20821 10625 20855 10659
rect 21189 10625 21223 10659
rect 21281 10625 21315 10659
rect 7757 10557 7791 10591
rect 8677 10557 8711 10591
rect 13737 10557 13771 10591
rect 14013 10557 14047 10591
rect 20729 10557 20763 10591
rect 16681 10489 16715 10523
rect 10517 10421 10551 10455
rect 11897 10421 11931 10455
rect 17141 10421 17175 10455
rect 21649 10421 21683 10455
rect 6469 10217 6503 10251
rect 10057 10217 10091 10251
rect 10333 10217 10367 10251
rect 14565 10217 14599 10251
rect 15945 10217 15979 10251
rect 18981 10217 19015 10251
rect 20361 10217 20395 10251
rect 21097 10217 21131 10251
rect 21465 10217 21499 10251
rect 9045 10149 9079 10183
rect 13461 10149 13495 10183
rect 13921 10149 13955 10183
rect 15577 10149 15611 10183
rect 19533 10149 19567 10183
rect 6745 10081 6779 10115
rect 11161 10081 11195 10115
rect 19625 10081 19659 10115
rect 9873 10013 9907 10047
rect 10885 10013 10919 10047
rect 13737 10013 13771 10047
rect 16589 10013 16623 10047
rect 16681 10013 16715 10047
rect 17141 10013 17175 10047
rect 17325 10013 17359 10047
rect 19404 10013 19438 10047
rect 22017 10013 22051 10047
rect 7021 9945 7055 9979
rect 8769 9945 8803 9979
rect 12909 9945 12943 9979
rect 18245 9945 18279 9979
rect 19257 9945 19291 9979
rect 19993 9945 20027 9979
rect 22293 9945 22327 9979
rect 24041 9945 24075 9979
rect 14289 9877 14323 9911
rect 17601 9877 17635 9911
rect 18613 9877 18647 9911
rect 7389 9673 7423 9707
rect 9781 9673 9815 9707
rect 11713 9673 11747 9707
rect 13645 9673 13679 9707
rect 14473 9673 14507 9707
rect 15301 9673 15335 9707
rect 17601 9673 17635 9707
rect 21189 9673 21223 9707
rect 22385 9673 22419 9707
rect 22753 9673 22787 9707
rect 7757 9605 7791 9639
rect 11069 9605 11103 9639
rect 15669 9605 15703 9639
rect 20177 9605 20211 9639
rect 20545 9605 20579 9639
rect 8217 9537 8251 9571
rect 8493 9537 8527 9571
rect 8585 9537 8619 9571
rect 10517 9537 10551 9571
rect 10701 9537 10735 9571
rect 12633 9537 12667 9571
rect 14473 9537 14507 9571
rect 16037 9537 16071 9571
rect 16681 9537 16715 9571
rect 19349 9537 19383 9571
rect 19717 9537 19751 9571
rect 19809 9537 19843 9571
rect 21005 9537 21039 9571
rect 23121 9537 23155 9571
rect 9045 9469 9079 9503
rect 9137 9469 9171 9503
rect 6469 9401 6503 9435
rect 11437 9401 11471 9435
rect 16865 9401 16899 9435
rect 19165 9401 19199 9435
rect 21557 9401 21591 9435
rect 7113 9333 7147 9367
rect 10057 9333 10091 9367
rect 12817 9333 12851 9367
rect 16405 9333 16439 9367
rect 17141 9333 17175 9367
rect 18613 9333 18647 9367
rect 22017 9333 22051 9367
rect 7389 9129 7423 9163
rect 8493 9129 8527 9163
rect 9045 9129 9079 9163
rect 10977 9129 11011 9163
rect 13829 9129 13863 9163
rect 14473 9129 14507 9163
rect 16313 9129 16347 9163
rect 19533 9129 19567 9163
rect 20177 9129 20211 9163
rect 22293 9129 22327 9163
rect 6929 9061 6963 9095
rect 11253 9061 11287 9095
rect 6561 8993 6595 9027
rect 10425 8993 10459 9027
rect 17417 8993 17451 9027
rect 19165 8993 19199 9027
rect 21097 8993 21131 9027
rect 7205 8925 7239 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 10057 8925 10091 8959
rect 12081 8925 12115 8959
rect 13645 8925 13679 8959
rect 14105 8925 14139 8959
rect 15485 8925 15519 8959
rect 15577 8925 15611 8959
rect 17141 8925 17175 8959
rect 21281 8925 21315 8959
rect 21833 8925 21867 8959
rect 22017 8925 22051 8959
rect 7849 8857 7883 8891
rect 9873 8857 9907 8891
rect 12725 8857 12759 8891
rect 16037 8857 16071 8891
rect 6193 8789 6227 8823
rect 13001 8789 13035 8823
rect 14933 8789 14967 8823
rect 16681 8789 16715 8823
rect 19901 8789 19935 8823
rect 8217 8585 8251 8619
rect 15669 8585 15703 8619
rect 17417 8585 17451 8619
rect 21741 8585 21775 8619
rect 22109 8585 22143 8619
rect 22845 8585 22879 8619
rect 9137 8517 9171 8551
rect 10701 8517 10735 8551
rect 21373 8517 21407 8551
rect 8585 8449 8619 8483
rect 8769 8449 8803 8483
rect 9965 8449 9999 8483
rect 10057 8449 10091 8483
rect 10241 8449 10275 8483
rect 10977 8449 11011 8483
rect 13001 8449 13035 8483
rect 16497 8449 16531 8483
rect 17141 8449 17175 8483
rect 18245 8449 18279 8483
rect 18429 8449 18463 8483
rect 19625 8449 19659 8483
rect 19717 8449 19751 8483
rect 19901 8449 19935 8483
rect 20269 8449 20303 8483
rect 20462 8449 20496 8483
rect 13277 8381 13311 8415
rect 15025 8381 15059 8415
rect 20821 8381 20855 8415
rect 7205 8245 7239 8279
rect 7941 8245 7975 8279
rect 9689 8245 9723 8279
rect 11989 8245 12023 8279
rect 12725 8245 12759 8279
rect 15301 8245 15335 8279
rect 16129 8245 16163 8279
rect 18521 8245 18555 8279
rect 19165 8245 19199 8279
rect 22477 8245 22511 8279
rect 7481 8041 7515 8075
rect 10057 8041 10091 8075
rect 11713 8041 11747 8075
rect 12265 8041 12299 8075
rect 14933 8041 14967 8075
rect 17509 8041 17543 8075
rect 18245 8041 18279 8075
rect 18870 8041 18904 8075
rect 19349 8041 19383 8075
rect 20453 8041 20487 8075
rect 21373 8041 21407 8075
rect 12541 7973 12575 8007
rect 18981 7973 19015 8007
rect 7113 7905 7147 7939
rect 13001 7905 13035 7939
rect 13277 7905 13311 7939
rect 15485 7905 15519 7939
rect 15945 7905 15979 7939
rect 19073 7905 19107 7939
rect 8309 7837 8343 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 11253 7837 11287 7871
rect 13829 7837 13863 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 16037 7837 16071 7871
rect 16497 7837 16531 7871
rect 16589 7837 16623 7871
rect 18705 7837 18739 7871
rect 21557 7837 21591 7871
rect 21741 7837 21775 7871
rect 22109 7837 22143 7871
rect 22201 7837 22235 7871
rect 7757 7769 7791 7803
rect 10701 7769 10735 7803
rect 17141 7769 17175 7803
rect 20085 7769 20119 7803
rect 9137 7701 9171 7735
rect 10333 7701 10367 7735
rect 17877 7701 17911 7735
rect 19717 7701 19751 7735
rect 8677 7497 8711 7531
rect 8953 7497 8987 7531
rect 10793 7497 10827 7531
rect 13553 7497 13587 7531
rect 14289 7497 14323 7531
rect 16129 7497 16163 7531
rect 17141 7497 17175 7531
rect 18337 7497 18371 7531
rect 19717 7497 19751 7531
rect 22753 7497 22787 7531
rect 10149 7429 10183 7463
rect 14841 7429 14875 7463
rect 15117 7429 15151 7463
rect 17417 7429 17451 7463
rect 19441 7429 19475 7463
rect 21833 7429 21867 7463
rect 7573 7361 7607 7395
rect 8309 7361 8343 7395
rect 9505 7361 9539 7395
rect 12725 7361 12759 7395
rect 13829 7361 13863 7395
rect 15577 7361 15611 7395
rect 16957 7361 16991 7395
rect 19165 7361 19199 7395
rect 20913 7361 20947 7395
rect 21281 7361 21315 7395
rect 21465 7361 21499 7395
rect 22293 7361 22327 7395
rect 7297 7293 7331 7327
rect 11069 7293 11103 7327
rect 12633 7293 12667 7327
rect 20821 7293 20855 7327
rect 11713 7225 11747 7259
rect 7665 7157 7699 7191
rect 12081 7157 12115 7191
rect 12909 7157 12943 7191
rect 14013 7157 14047 7191
rect 16497 7157 16531 7191
rect 20545 7157 20579 7191
rect 22477 7157 22511 7191
rect 14657 6953 14691 6987
rect 17049 6953 17083 6987
rect 17509 6953 17543 6987
rect 20453 6953 20487 6987
rect 15577 6885 15611 6919
rect 18429 6885 18463 6919
rect 6653 6817 6687 6851
rect 12081 6817 12115 6851
rect 14381 6817 14415 6851
rect 16037 6817 16071 6851
rect 16589 6817 16623 6851
rect 19257 6817 19291 6851
rect 19717 6817 19751 6851
rect 21465 6817 21499 6851
rect 23213 6817 23247 6851
rect 23489 6817 23523 6851
rect 7757 6749 7791 6783
rect 7941 6749 7975 6783
rect 8125 6749 8159 6783
rect 8585 6749 8619 6783
rect 8677 6749 8711 6783
rect 10517 6749 10551 6783
rect 12357 6749 12391 6783
rect 16129 6749 16163 6783
rect 17785 6749 17819 6783
rect 19441 6749 19475 6783
rect 19809 6749 19843 6783
rect 21189 6749 21223 6783
rect 7297 6681 7331 6715
rect 10057 6681 10091 6715
rect 12633 6681 12667 6715
rect 7021 6613 7055 6647
rect 9229 6613 9263 6647
rect 11161 6613 11195 6647
rect 11713 6613 11747 6647
rect 17969 6613 18003 6647
rect 19073 6613 19107 6647
rect 5917 6409 5951 6443
rect 9689 6409 9723 6443
rect 11713 6409 11747 6443
rect 14841 6409 14875 6443
rect 17693 6409 17727 6443
rect 22661 6409 22695 6443
rect 11345 6341 11379 6375
rect 17141 6341 17175 6375
rect 19073 6341 19107 6375
rect 21649 6341 21683 6375
rect 5733 6273 5767 6307
rect 9965 6273 9999 6307
rect 10793 6273 10827 6307
rect 13093 6273 13127 6307
rect 13461 6273 13495 6307
rect 14657 6273 14691 6307
rect 16313 6273 16347 6307
rect 16681 6273 16715 6307
rect 21741 6273 21775 6307
rect 7113 6205 7147 6239
rect 7389 6205 7423 6239
rect 9137 6205 9171 6239
rect 10517 6205 10551 6239
rect 10977 6205 11011 6239
rect 12633 6205 12667 6239
rect 13553 6205 13587 6239
rect 16405 6205 16439 6239
rect 16773 6205 16807 6239
rect 18797 6205 18831 6239
rect 20821 6205 20855 6239
rect 15393 6137 15427 6171
rect 6469 6069 6503 6103
rect 11989 6069 12023 6103
rect 13921 6069 13955 6103
rect 14381 6069 14415 6103
rect 15761 6069 15795 6103
rect 18245 6069 18279 6103
rect 21189 6069 21223 6103
rect 5733 5865 5767 5899
rect 6469 5865 6503 5899
rect 6837 5865 6871 5899
rect 8033 5865 8067 5899
rect 8677 5865 8711 5899
rect 10149 5865 10183 5899
rect 12449 5865 12483 5899
rect 14289 5865 14323 5899
rect 15761 5865 15795 5899
rect 18245 5865 18279 5899
rect 19809 5865 19843 5899
rect 20361 5865 20395 5899
rect 21189 5865 21223 5899
rect 21649 5865 21683 5899
rect 9321 5797 9355 5831
rect 14933 5797 14967 5831
rect 10793 5729 10827 5763
rect 11345 5729 11379 5763
rect 12081 5729 12115 5763
rect 18889 5729 18923 5763
rect 19441 5729 19475 5763
rect 7941 5661 7975 5695
rect 10057 5661 10091 5695
rect 11529 5661 11563 5695
rect 12909 5661 12943 5695
rect 13001 5661 13035 5695
rect 13185 5661 13219 5695
rect 15577 5661 15611 5695
rect 17141 5661 17175 5695
rect 17417 5661 17451 5695
rect 17601 5661 17635 5695
rect 18981 5661 19015 5695
rect 7757 5593 7791 5627
rect 9873 5593 9907 5627
rect 11621 5593 11655 5627
rect 11713 5593 11747 5627
rect 13645 5593 13679 5627
rect 16589 5593 16623 5627
rect 7205 5525 7239 5559
rect 14013 5525 14047 5559
rect 16037 5525 16071 5559
rect 18521 5525 18555 5559
rect 21925 5525 21959 5559
rect 22293 5525 22327 5559
rect 7205 5321 7239 5355
rect 7757 5321 7791 5355
rect 8217 5321 8251 5355
rect 9045 5321 9079 5355
rect 9873 5321 9907 5355
rect 11805 5321 11839 5355
rect 14197 5321 14231 5355
rect 14749 5321 14783 5355
rect 17417 5321 17451 5355
rect 19257 5321 19291 5355
rect 20637 5321 20671 5355
rect 20913 5321 20947 5355
rect 21741 5321 21775 5355
rect 15761 5253 15795 5287
rect 16313 5253 16347 5287
rect 20269 5253 20303 5287
rect 9321 5185 9355 5219
rect 10333 5185 10367 5219
rect 10793 5185 10827 5219
rect 10977 5185 11011 5219
rect 11345 5185 11379 5219
rect 12725 5185 12759 5219
rect 14013 5185 14047 5219
rect 15117 5185 15151 5219
rect 16681 5185 16715 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 19809 5185 19843 5219
rect 11253 5117 11287 5151
rect 12633 5117 12667 5151
rect 16589 5117 16623 5151
rect 18337 5117 18371 5151
rect 18705 5117 18739 5151
rect 19717 5117 19751 5151
rect 21281 5117 21315 5151
rect 8677 4981 8711 5015
rect 9505 4981 9539 5015
rect 13645 4981 13679 5015
rect 16865 4981 16899 5015
rect 7849 4777 7883 4811
rect 8953 4777 8987 4811
rect 12633 4777 12667 4811
rect 13369 4777 13403 4811
rect 14565 4777 14599 4811
rect 18153 4777 18187 4811
rect 19165 4777 19199 4811
rect 19901 4777 19935 4811
rect 20177 4777 20211 4811
rect 8585 4709 8619 4743
rect 8217 4641 8251 4675
rect 11529 4641 11563 4675
rect 15485 4641 15519 4675
rect 16129 4641 16163 4675
rect 17877 4641 17911 4675
rect 21097 4641 21131 4675
rect 21465 4641 21499 4675
rect 10241 4573 10275 4607
rect 11069 4573 11103 4607
rect 11345 4573 11379 4607
rect 13001 4573 13035 4607
rect 15853 4573 15887 4607
rect 18705 4573 18739 4607
rect 19717 4573 19751 4607
rect 10517 4505 10551 4539
rect 14933 4505 14967 4539
rect 9229 4437 9263 4471
rect 11805 4437 11839 4471
rect 14105 4437 14139 4471
rect 18889 4437 18923 4471
rect 7849 4233 7883 4267
rect 15577 4233 15611 4267
rect 17417 4233 17451 4267
rect 19349 4233 19383 4267
rect 20453 4233 20487 4267
rect 9137 4165 9171 4199
rect 11529 4165 11563 4199
rect 16405 4165 16439 4199
rect 8125 4097 8159 4131
rect 8309 4097 8343 4131
rect 11897 4097 11931 4131
rect 14013 4097 14047 4131
rect 15393 4097 15427 4131
rect 17049 4097 17083 4131
rect 18705 4097 18739 4131
rect 19625 4097 19659 4131
rect 20085 4097 20119 4131
rect 7481 4029 7515 4063
rect 8677 4029 8711 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 18245 4029 18279 4063
rect 15117 3961 15151 3995
rect 19809 3961 19843 3995
rect 12909 3893 12943 3927
rect 13645 3893 13679 3927
rect 14473 3893 14507 3927
rect 15945 3893 15979 3927
rect 8585 3689 8619 3723
rect 12725 3689 12759 3723
rect 14473 3689 14507 3723
rect 15945 3689 15979 3723
rect 18797 3689 18831 3723
rect 8217 3621 8251 3655
rect 15577 3621 15611 3655
rect 14105 3553 14139 3587
rect 16773 3553 16807 3587
rect 18153 3553 18187 3587
rect 19165 3553 19199 3587
rect 10149 3485 10183 3519
rect 13093 3485 13127 3519
rect 13645 3485 13679 3519
rect 16405 3485 16439 3519
rect 19625 3485 19659 3519
rect 8953 3417 8987 3451
rect 10425 3417 10459 3451
rect 12173 3417 12207 3451
rect 9229 3349 9263 3383
rect 13185 3349 13219 3383
rect 14933 3349 14967 3383
rect 8861 3145 8895 3179
rect 10977 3145 11011 3179
rect 12817 3145 12851 3179
rect 17417 3145 17451 3179
rect 19073 3145 19107 3179
rect 19441 3145 19475 3179
rect 9781 3077 9815 3111
rect 14013 3077 14047 3111
rect 9689 3009 9723 3043
rect 10517 3009 10551 3043
rect 10609 3009 10643 3043
rect 12541 3009 12575 3043
rect 12633 3009 12667 3043
rect 16681 3009 16715 3043
rect 18245 3009 18279 3043
rect 11437 2941 11471 2975
rect 13737 2941 13771 2975
rect 15761 2941 15795 2975
rect 16589 2941 16623 2975
rect 18705 2941 18739 2975
rect 11989 2873 12023 2907
rect 12541 2873 12575 2907
rect 13185 2873 13219 2907
rect 18429 2873 18463 2907
rect 9321 2805 9355 2839
rect 16221 2805 16255 2839
rect 16865 2805 16899 2839
rect 8953 2601 8987 2635
rect 10149 2601 10183 2635
rect 13185 2601 13219 2635
rect 14289 2601 14323 2635
rect 14841 2601 14875 2635
rect 16037 2601 16071 2635
rect 18705 2601 18739 2635
rect 10425 2533 10459 2567
rect 12265 2533 12299 2567
rect 13967 2533 14001 2567
rect 14105 2533 14139 2567
rect 19717 2533 19751 2567
rect 7941 2465 7975 2499
rect 11069 2465 11103 2499
rect 11437 2465 11471 2499
rect 14197 2465 14231 2499
rect 17785 2465 17819 2499
rect 8677 2397 8711 2431
rect 9965 2397 9999 2431
rect 10977 2397 11011 2431
rect 11253 2397 11287 2431
rect 13461 2397 13495 2431
rect 16405 2397 16439 2431
rect 17325 2397 17359 2431
rect 18521 2397 18555 2431
rect 19349 2397 19383 2431
rect 9413 2329 9447 2363
rect 13829 2329 13863 2363
rect 16681 2329 16715 2363
rect 18981 2329 19015 2363
rect 8309 2261 8343 2295
rect 20085 2261 20119 2295
<< metal1 >>
rect 1104 29402 28336 29424
rect 1104 29350 1782 29402
rect 1834 29350 1846 29402
rect 1898 29350 1910 29402
rect 1962 29350 1974 29402
rect 2026 29350 4782 29402
rect 4834 29350 4846 29402
rect 4898 29350 4910 29402
rect 4962 29350 4974 29402
rect 5026 29350 7782 29402
rect 7834 29350 7846 29402
rect 7898 29350 7910 29402
rect 7962 29350 7974 29402
rect 8026 29350 10782 29402
rect 10834 29350 10846 29402
rect 10898 29350 10910 29402
rect 10962 29350 10974 29402
rect 11026 29350 13782 29402
rect 13834 29350 13846 29402
rect 13898 29350 13910 29402
rect 13962 29350 13974 29402
rect 14026 29350 16782 29402
rect 16834 29350 16846 29402
rect 16898 29350 16910 29402
rect 16962 29350 16974 29402
rect 17026 29350 19782 29402
rect 19834 29350 19846 29402
rect 19898 29350 19910 29402
rect 19962 29350 19974 29402
rect 20026 29350 22782 29402
rect 22834 29350 22846 29402
rect 22898 29350 22910 29402
rect 22962 29350 22974 29402
rect 23026 29350 25782 29402
rect 25834 29350 25846 29402
rect 25898 29350 25910 29402
rect 25962 29350 25974 29402
rect 26026 29350 28336 29402
rect 1104 29328 28336 29350
rect 1104 28858 28336 28880
rect 1104 28806 3282 28858
rect 3334 28806 3346 28858
rect 3398 28806 3410 28858
rect 3462 28806 3474 28858
rect 3526 28806 6282 28858
rect 6334 28806 6346 28858
rect 6398 28806 6410 28858
rect 6462 28806 6474 28858
rect 6526 28806 9282 28858
rect 9334 28806 9346 28858
rect 9398 28806 9410 28858
rect 9462 28806 9474 28858
rect 9526 28806 12282 28858
rect 12334 28806 12346 28858
rect 12398 28806 12410 28858
rect 12462 28806 12474 28858
rect 12526 28806 15282 28858
rect 15334 28806 15346 28858
rect 15398 28806 15410 28858
rect 15462 28806 15474 28858
rect 15526 28806 18282 28858
rect 18334 28806 18346 28858
rect 18398 28806 18410 28858
rect 18462 28806 18474 28858
rect 18526 28806 21282 28858
rect 21334 28806 21346 28858
rect 21398 28806 21410 28858
rect 21462 28806 21474 28858
rect 21526 28806 24282 28858
rect 24334 28806 24346 28858
rect 24398 28806 24410 28858
rect 24462 28806 24474 28858
rect 24526 28806 27282 28858
rect 27334 28806 27346 28858
rect 27398 28806 27410 28858
rect 27462 28806 27474 28858
rect 27526 28806 28336 28858
rect 1104 28784 28336 28806
rect 1104 28314 28336 28336
rect 1104 28262 1782 28314
rect 1834 28262 1846 28314
rect 1898 28262 1910 28314
rect 1962 28262 1974 28314
rect 2026 28262 4782 28314
rect 4834 28262 4846 28314
rect 4898 28262 4910 28314
rect 4962 28262 4974 28314
rect 5026 28262 7782 28314
rect 7834 28262 7846 28314
rect 7898 28262 7910 28314
rect 7962 28262 7974 28314
rect 8026 28262 10782 28314
rect 10834 28262 10846 28314
rect 10898 28262 10910 28314
rect 10962 28262 10974 28314
rect 11026 28262 13782 28314
rect 13834 28262 13846 28314
rect 13898 28262 13910 28314
rect 13962 28262 13974 28314
rect 14026 28262 16782 28314
rect 16834 28262 16846 28314
rect 16898 28262 16910 28314
rect 16962 28262 16974 28314
rect 17026 28262 19782 28314
rect 19834 28262 19846 28314
rect 19898 28262 19910 28314
rect 19962 28262 19974 28314
rect 20026 28262 22782 28314
rect 22834 28262 22846 28314
rect 22898 28262 22910 28314
rect 22962 28262 22974 28314
rect 23026 28262 25782 28314
rect 25834 28262 25846 28314
rect 25898 28262 25910 28314
rect 25962 28262 25974 28314
rect 26026 28262 28336 28314
rect 1104 28240 28336 28262
rect 1104 27770 28336 27792
rect 1104 27718 3282 27770
rect 3334 27718 3346 27770
rect 3398 27718 3410 27770
rect 3462 27718 3474 27770
rect 3526 27718 6282 27770
rect 6334 27718 6346 27770
rect 6398 27718 6410 27770
rect 6462 27718 6474 27770
rect 6526 27718 9282 27770
rect 9334 27718 9346 27770
rect 9398 27718 9410 27770
rect 9462 27718 9474 27770
rect 9526 27718 12282 27770
rect 12334 27718 12346 27770
rect 12398 27718 12410 27770
rect 12462 27718 12474 27770
rect 12526 27718 15282 27770
rect 15334 27718 15346 27770
rect 15398 27718 15410 27770
rect 15462 27718 15474 27770
rect 15526 27718 18282 27770
rect 18334 27718 18346 27770
rect 18398 27718 18410 27770
rect 18462 27718 18474 27770
rect 18526 27718 21282 27770
rect 21334 27718 21346 27770
rect 21398 27718 21410 27770
rect 21462 27718 21474 27770
rect 21526 27718 24282 27770
rect 24334 27718 24346 27770
rect 24398 27718 24410 27770
rect 24462 27718 24474 27770
rect 24526 27718 27282 27770
rect 27334 27718 27346 27770
rect 27398 27718 27410 27770
rect 27462 27718 27474 27770
rect 27526 27718 28336 27770
rect 1104 27696 28336 27718
rect 23198 27412 23204 27464
rect 23256 27452 23262 27464
rect 23753 27455 23811 27461
rect 23753 27452 23765 27455
rect 23256 27424 23765 27452
rect 23256 27412 23262 27424
rect 23753 27421 23765 27424
rect 23799 27452 23811 27455
rect 24578 27452 24584 27464
rect 23799 27424 24584 27452
rect 23799 27421 23811 27424
rect 23753 27415 23811 27421
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 23106 27384 23112 27396
rect 23067 27356 23112 27384
rect 23106 27344 23112 27356
rect 23164 27344 23170 27396
rect 1104 27226 28336 27248
rect 1104 27174 1782 27226
rect 1834 27174 1846 27226
rect 1898 27174 1910 27226
rect 1962 27174 1974 27226
rect 2026 27174 4782 27226
rect 4834 27174 4846 27226
rect 4898 27174 4910 27226
rect 4962 27174 4974 27226
rect 5026 27174 7782 27226
rect 7834 27174 7846 27226
rect 7898 27174 7910 27226
rect 7962 27174 7974 27226
rect 8026 27174 10782 27226
rect 10834 27174 10846 27226
rect 10898 27174 10910 27226
rect 10962 27174 10974 27226
rect 11026 27174 13782 27226
rect 13834 27174 13846 27226
rect 13898 27174 13910 27226
rect 13962 27174 13974 27226
rect 14026 27174 16782 27226
rect 16834 27174 16846 27226
rect 16898 27174 16910 27226
rect 16962 27174 16974 27226
rect 17026 27174 19782 27226
rect 19834 27174 19846 27226
rect 19898 27174 19910 27226
rect 19962 27174 19974 27226
rect 20026 27174 22782 27226
rect 22834 27174 22846 27226
rect 22898 27174 22910 27226
rect 22962 27174 22974 27226
rect 23026 27174 25782 27226
rect 25834 27174 25846 27226
rect 25898 27174 25910 27226
rect 25962 27174 25974 27226
rect 26026 27174 28336 27226
rect 1104 27152 28336 27174
rect 23198 27112 23204 27124
rect 23159 27084 23204 27112
rect 23198 27072 23204 27084
rect 23256 27072 23262 27124
rect 1104 26682 28336 26704
rect 1104 26630 3282 26682
rect 3334 26630 3346 26682
rect 3398 26630 3410 26682
rect 3462 26630 3474 26682
rect 3526 26630 6282 26682
rect 6334 26630 6346 26682
rect 6398 26630 6410 26682
rect 6462 26630 6474 26682
rect 6526 26630 9282 26682
rect 9334 26630 9346 26682
rect 9398 26630 9410 26682
rect 9462 26630 9474 26682
rect 9526 26630 12282 26682
rect 12334 26630 12346 26682
rect 12398 26630 12410 26682
rect 12462 26630 12474 26682
rect 12526 26630 15282 26682
rect 15334 26630 15346 26682
rect 15398 26630 15410 26682
rect 15462 26630 15474 26682
rect 15526 26630 18282 26682
rect 18334 26630 18346 26682
rect 18398 26630 18410 26682
rect 18462 26630 18474 26682
rect 18526 26630 21282 26682
rect 21334 26630 21346 26682
rect 21398 26630 21410 26682
rect 21462 26630 21474 26682
rect 21526 26630 24282 26682
rect 24334 26630 24346 26682
rect 24398 26630 24410 26682
rect 24462 26630 24474 26682
rect 24526 26630 27282 26682
rect 27334 26630 27346 26682
rect 27398 26630 27410 26682
rect 27462 26630 27474 26682
rect 27526 26630 28336 26682
rect 1104 26608 28336 26630
rect 1104 26138 28336 26160
rect 1104 26086 1782 26138
rect 1834 26086 1846 26138
rect 1898 26086 1910 26138
rect 1962 26086 1974 26138
rect 2026 26086 4782 26138
rect 4834 26086 4846 26138
rect 4898 26086 4910 26138
rect 4962 26086 4974 26138
rect 5026 26086 7782 26138
rect 7834 26086 7846 26138
rect 7898 26086 7910 26138
rect 7962 26086 7974 26138
rect 8026 26086 10782 26138
rect 10834 26086 10846 26138
rect 10898 26086 10910 26138
rect 10962 26086 10974 26138
rect 11026 26086 13782 26138
rect 13834 26086 13846 26138
rect 13898 26086 13910 26138
rect 13962 26086 13974 26138
rect 14026 26086 16782 26138
rect 16834 26086 16846 26138
rect 16898 26086 16910 26138
rect 16962 26086 16974 26138
rect 17026 26086 19782 26138
rect 19834 26086 19846 26138
rect 19898 26086 19910 26138
rect 19962 26086 19974 26138
rect 20026 26086 22782 26138
rect 22834 26086 22846 26138
rect 22898 26086 22910 26138
rect 22962 26086 22974 26138
rect 23026 26086 25782 26138
rect 25834 26086 25846 26138
rect 25898 26086 25910 26138
rect 25962 26086 25974 26138
rect 26026 26086 28336 26138
rect 1104 26064 28336 26086
rect 1104 25594 28336 25616
rect 1104 25542 3282 25594
rect 3334 25542 3346 25594
rect 3398 25542 3410 25594
rect 3462 25542 3474 25594
rect 3526 25542 6282 25594
rect 6334 25542 6346 25594
rect 6398 25542 6410 25594
rect 6462 25542 6474 25594
rect 6526 25542 9282 25594
rect 9334 25542 9346 25594
rect 9398 25542 9410 25594
rect 9462 25542 9474 25594
rect 9526 25542 12282 25594
rect 12334 25542 12346 25594
rect 12398 25542 12410 25594
rect 12462 25542 12474 25594
rect 12526 25542 15282 25594
rect 15334 25542 15346 25594
rect 15398 25542 15410 25594
rect 15462 25542 15474 25594
rect 15526 25542 18282 25594
rect 18334 25542 18346 25594
rect 18398 25542 18410 25594
rect 18462 25542 18474 25594
rect 18526 25542 21282 25594
rect 21334 25542 21346 25594
rect 21398 25542 21410 25594
rect 21462 25542 21474 25594
rect 21526 25542 24282 25594
rect 24334 25542 24346 25594
rect 24398 25542 24410 25594
rect 24462 25542 24474 25594
rect 24526 25542 27282 25594
rect 27334 25542 27346 25594
rect 27398 25542 27410 25594
rect 27462 25542 27474 25594
rect 27526 25542 28336 25594
rect 1104 25520 28336 25542
rect 1104 25050 28336 25072
rect 1104 24998 1782 25050
rect 1834 24998 1846 25050
rect 1898 24998 1910 25050
rect 1962 24998 1974 25050
rect 2026 24998 4782 25050
rect 4834 24998 4846 25050
rect 4898 24998 4910 25050
rect 4962 24998 4974 25050
rect 5026 24998 7782 25050
rect 7834 24998 7846 25050
rect 7898 24998 7910 25050
rect 7962 24998 7974 25050
rect 8026 24998 10782 25050
rect 10834 24998 10846 25050
rect 10898 24998 10910 25050
rect 10962 24998 10974 25050
rect 11026 24998 13782 25050
rect 13834 24998 13846 25050
rect 13898 24998 13910 25050
rect 13962 24998 13974 25050
rect 14026 24998 16782 25050
rect 16834 24998 16846 25050
rect 16898 24998 16910 25050
rect 16962 24998 16974 25050
rect 17026 24998 19782 25050
rect 19834 24998 19846 25050
rect 19898 24998 19910 25050
rect 19962 24998 19974 25050
rect 20026 24998 22782 25050
rect 22834 24998 22846 25050
rect 22898 24998 22910 25050
rect 22962 24998 22974 25050
rect 23026 24998 25782 25050
rect 25834 24998 25846 25050
rect 25898 24998 25910 25050
rect 25962 24998 25974 25050
rect 26026 24998 28336 25050
rect 1104 24976 28336 24998
rect 1104 24506 28336 24528
rect 1104 24454 3282 24506
rect 3334 24454 3346 24506
rect 3398 24454 3410 24506
rect 3462 24454 3474 24506
rect 3526 24454 6282 24506
rect 6334 24454 6346 24506
rect 6398 24454 6410 24506
rect 6462 24454 6474 24506
rect 6526 24454 9282 24506
rect 9334 24454 9346 24506
rect 9398 24454 9410 24506
rect 9462 24454 9474 24506
rect 9526 24454 12282 24506
rect 12334 24454 12346 24506
rect 12398 24454 12410 24506
rect 12462 24454 12474 24506
rect 12526 24454 15282 24506
rect 15334 24454 15346 24506
rect 15398 24454 15410 24506
rect 15462 24454 15474 24506
rect 15526 24454 18282 24506
rect 18334 24454 18346 24506
rect 18398 24454 18410 24506
rect 18462 24454 18474 24506
rect 18526 24454 21282 24506
rect 21334 24454 21346 24506
rect 21398 24454 21410 24506
rect 21462 24454 21474 24506
rect 21526 24454 24282 24506
rect 24334 24454 24346 24506
rect 24398 24454 24410 24506
rect 24462 24454 24474 24506
rect 24526 24454 27282 24506
rect 27334 24454 27346 24506
rect 27398 24454 27410 24506
rect 27462 24454 27474 24506
rect 27526 24454 28336 24506
rect 1104 24432 28336 24454
rect 1104 23962 28336 23984
rect 1104 23910 1782 23962
rect 1834 23910 1846 23962
rect 1898 23910 1910 23962
rect 1962 23910 1974 23962
rect 2026 23910 4782 23962
rect 4834 23910 4846 23962
rect 4898 23910 4910 23962
rect 4962 23910 4974 23962
rect 5026 23910 7782 23962
rect 7834 23910 7846 23962
rect 7898 23910 7910 23962
rect 7962 23910 7974 23962
rect 8026 23910 10782 23962
rect 10834 23910 10846 23962
rect 10898 23910 10910 23962
rect 10962 23910 10974 23962
rect 11026 23910 13782 23962
rect 13834 23910 13846 23962
rect 13898 23910 13910 23962
rect 13962 23910 13974 23962
rect 14026 23910 16782 23962
rect 16834 23910 16846 23962
rect 16898 23910 16910 23962
rect 16962 23910 16974 23962
rect 17026 23910 19782 23962
rect 19834 23910 19846 23962
rect 19898 23910 19910 23962
rect 19962 23910 19974 23962
rect 20026 23910 22782 23962
rect 22834 23910 22846 23962
rect 22898 23910 22910 23962
rect 22962 23910 22974 23962
rect 23026 23910 25782 23962
rect 25834 23910 25846 23962
rect 25898 23910 25910 23962
rect 25962 23910 25974 23962
rect 26026 23910 28336 23962
rect 1104 23888 28336 23910
rect 1104 23418 28336 23440
rect 1104 23366 3282 23418
rect 3334 23366 3346 23418
rect 3398 23366 3410 23418
rect 3462 23366 3474 23418
rect 3526 23366 6282 23418
rect 6334 23366 6346 23418
rect 6398 23366 6410 23418
rect 6462 23366 6474 23418
rect 6526 23366 9282 23418
rect 9334 23366 9346 23418
rect 9398 23366 9410 23418
rect 9462 23366 9474 23418
rect 9526 23366 12282 23418
rect 12334 23366 12346 23418
rect 12398 23366 12410 23418
rect 12462 23366 12474 23418
rect 12526 23366 15282 23418
rect 15334 23366 15346 23418
rect 15398 23366 15410 23418
rect 15462 23366 15474 23418
rect 15526 23366 18282 23418
rect 18334 23366 18346 23418
rect 18398 23366 18410 23418
rect 18462 23366 18474 23418
rect 18526 23366 21282 23418
rect 21334 23366 21346 23418
rect 21398 23366 21410 23418
rect 21462 23366 21474 23418
rect 21526 23366 24282 23418
rect 24334 23366 24346 23418
rect 24398 23366 24410 23418
rect 24462 23366 24474 23418
rect 24526 23366 27282 23418
rect 27334 23366 27346 23418
rect 27398 23366 27410 23418
rect 27462 23366 27474 23418
rect 27526 23366 28336 23418
rect 1104 23344 28336 23366
rect 1104 22874 28336 22896
rect 1104 22822 1782 22874
rect 1834 22822 1846 22874
rect 1898 22822 1910 22874
rect 1962 22822 1974 22874
rect 2026 22822 4782 22874
rect 4834 22822 4846 22874
rect 4898 22822 4910 22874
rect 4962 22822 4974 22874
rect 5026 22822 7782 22874
rect 7834 22822 7846 22874
rect 7898 22822 7910 22874
rect 7962 22822 7974 22874
rect 8026 22822 10782 22874
rect 10834 22822 10846 22874
rect 10898 22822 10910 22874
rect 10962 22822 10974 22874
rect 11026 22822 13782 22874
rect 13834 22822 13846 22874
rect 13898 22822 13910 22874
rect 13962 22822 13974 22874
rect 14026 22822 16782 22874
rect 16834 22822 16846 22874
rect 16898 22822 16910 22874
rect 16962 22822 16974 22874
rect 17026 22822 19782 22874
rect 19834 22822 19846 22874
rect 19898 22822 19910 22874
rect 19962 22822 19974 22874
rect 20026 22822 22782 22874
rect 22834 22822 22846 22874
rect 22898 22822 22910 22874
rect 22962 22822 22974 22874
rect 23026 22822 25782 22874
rect 25834 22822 25846 22874
rect 25898 22822 25910 22874
rect 25962 22822 25974 22874
rect 26026 22822 28336 22874
rect 1104 22800 28336 22822
rect 1104 22330 28336 22352
rect 1104 22278 3282 22330
rect 3334 22278 3346 22330
rect 3398 22278 3410 22330
rect 3462 22278 3474 22330
rect 3526 22278 6282 22330
rect 6334 22278 6346 22330
rect 6398 22278 6410 22330
rect 6462 22278 6474 22330
rect 6526 22278 9282 22330
rect 9334 22278 9346 22330
rect 9398 22278 9410 22330
rect 9462 22278 9474 22330
rect 9526 22278 12282 22330
rect 12334 22278 12346 22330
rect 12398 22278 12410 22330
rect 12462 22278 12474 22330
rect 12526 22278 15282 22330
rect 15334 22278 15346 22330
rect 15398 22278 15410 22330
rect 15462 22278 15474 22330
rect 15526 22278 18282 22330
rect 18334 22278 18346 22330
rect 18398 22278 18410 22330
rect 18462 22278 18474 22330
rect 18526 22278 21282 22330
rect 21334 22278 21346 22330
rect 21398 22278 21410 22330
rect 21462 22278 21474 22330
rect 21526 22278 24282 22330
rect 24334 22278 24346 22330
rect 24398 22278 24410 22330
rect 24462 22278 24474 22330
rect 24526 22278 27282 22330
rect 27334 22278 27346 22330
rect 27398 22278 27410 22330
rect 27462 22278 27474 22330
rect 27526 22278 28336 22330
rect 1104 22256 28336 22278
rect 1104 21786 28336 21808
rect 1104 21734 1782 21786
rect 1834 21734 1846 21786
rect 1898 21734 1910 21786
rect 1962 21734 1974 21786
rect 2026 21734 4782 21786
rect 4834 21734 4846 21786
rect 4898 21734 4910 21786
rect 4962 21734 4974 21786
rect 5026 21734 7782 21786
rect 7834 21734 7846 21786
rect 7898 21734 7910 21786
rect 7962 21734 7974 21786
rect 8026 21734 10782 21786
rect 10834 21734 10846 21786
rect 10898 21734 10910 21786
rect 10962 21734 10974 21786
rect 11026 21734 13782 21786
rect 13834 21734 13846 21786
rect 13898 21734 13910 21786
rect 13962 21734 13974 21786
rect 14026 21734 16782 21786
rect 16834 21734 16846 21786
rect 16898 21734 16910 21786
rect 16962 21734 16974 21786
rect 17026 21734 19782 21786
rect 19834 21734 19846 21786
rect 19898 21734 19910 21786
rect 19962 21734 19974 21786
rect 20026 21734 22782 21786
rect 22834 21734 22846 21786
rect 22898 21734 22910 21786
rect 22962 21734 22974 21786
rect 23026 21734 25782 21786
rect 25834 21734 25846 21786
rect 25898 21734 25910 21786
rect 25962 21734 25974 21786
rect 26026 21734 28336 21786
rect 1104 21712 28336 21734
rect 1104 21242 28336 21264
rect 1104 21190 3282 21242
rect 3334 21190 3346 21242
rect 3398 21190 3410 21242
rect 3462 21190 3474 21242
rect 3526 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 6410 21242
rect 6462 21190 6474 21242
rect 6526 21190 9282 21242
rect 9334 21190 9346 21242
rect 9398 21190 9410 21242
rect 9462 21190 9474 21242
rect 9526 21190 12282 21242
rect 12334 21190 12346 21242
rect 12398 21190 12410 21242
rect 12462 21190 12474 21242
rect 12526 21190 15282 21242
rect 15334 21190 15346 21242
rect 15398 21190 15410 21242
rect 15462 21190 15474 21242
rect 15526 21190 18282 21242
rect 18334 21190 18346 21242
rect 18398 21190 18410 21242
rect 18462 21190 18474 21242
rect 18526 21190 21282 21242
rect 21334 21190 21346 21242
rect 21398 21190 21410 21242
rect 21462 21190 21474 21242
rect 21526 21190 24282 21242
rect 24334 21190 24346 21242
rect 24398 21190 24410 21242
rect 24462 21190 24474 21242
rect 24526 21190 27282 21242
rect 27334 21190 27346 21242
rect 27398 21190 27410 21242
rect 27462 21190 27474 21242
rect 27526 21190 28336 21242
rect 1104 21168 28336 21190
rect 1104 20698 28336 20720
rect 1104 20646 1782 20698
rect 1834 20646 1846 20698
rect 1898 20646 1910 20698
rect 1962 20646 1974 20698
rect 2026 20646 4782 20698
rect 4834 20646 4846 20698
rect 4898 20646 4910 20698
rect 4962 20646 4974 20698
rect 5026 20646 7782 20698
rect 7834 20646 7846 20698
rect 7898 20646 7910 20698
rect 7962 20646 7974 20698
rect 8026 20646 10782 20698
rect 10834 20646 10846 20698
rect 10898 20646 10910 20698
rect 10962 20646 10974 20698
rect 11026 20646 13782 20698
rect 13834 20646 13846 20698
rect 13898 20646 13910 20698
rect 13962 20646 13974 20698
rect 14026 20646 16782 20698
rect 16834 20646 16846 20698
rect 16898 20646 16910 20698
rect 16962 20646 16974 20698
rect 17026 20646 19782 20698
rect 19834 20646 19846 20698
rect 19898 20646 19910 20698
rect 19962 20646 19974 20698
rect 20026 20646 22782 20698
rect 22834 20646 22846 20698
rect 22898 20646 22910 20698
rect 22962 20646 22974 20698
rect 23026 20646 25782 20698
rect 25834 20646 25846 20698
rect 25898 20646 25910 20698
rect 25962 20646 25974 20698
rect 26026 20646 28336 20698
rect 1104 20624 28336 20646
rect 1104 20154 28336 20176
rect 1104 20102 3282 20154
rect 3334 20102 3346 20154
rect 3398 20102 3410 20154
rect 3462 20102 3474 20154
rect 3526 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 6410 20154
rect 6462 20102 6474 20154
rect 6526 20102 9282 20154
rect 9334 20102 9346 20154
rect 9398 20102 9410 20154
rect 9462 20102 9474 20154
rect 9526 20102 12282 20154
rect 12334 20102 12346 20154
rect 12398 20102 12410 20154
rect 12462 20102 12474 20154
rect 12526 20102 15282 20154
rect 15334 20102 15346 20154
rect 15398 20102 15410 20154
rect 15462 20102 15474 20154
rect 15526 20102 18282 20154
rect 18334 20102 18346 20154
rect 18398 20102 18410 20154
rect 18462 20102 18474 20154
rect 18526 20102 21282 20154
rect 21334 20102 21346 20154
rect 21398 20102 21410 20154
rect 21462 20102 21474 20154
rect 21526 20102 24282 20154
rect 24334 20102 24346 20154
rect 24398 20102 24410 20154
rect 24462 20102 24474 20154
rect 24526 20102 27282 20154
rect 27334 20102 27346 20154
rect 27398 20102 27410 20154
rect 27462 20102 27474 20154
rect 27526 20102 28336 20154
rect 1104 20080 28336 20102
rect 1104 19610 28336 19632
rect 1104 19558 1782 19610
rect 1834 19558 1846 19610
rect 1898 19558 1910 19610
rect 1962 19558 1974 19610
rect 2026 19558 4782 19610
rect 4834 19558 4846 19610
rect 4898 19558 4910 19610
rect 4962 19558 4974 19610
rect 5026 19558 7782 19610
rect 7834 19558 7846 19610
rect 7898 19558 7910 19610
rect 7962 19558 7974 19610
rect 8026 19558 10782 19610
rect 10834 19558 10846 19610
rect 10898 19558 10910 19610
rect 10962 19558 10974 19610
rect 11026 19558 13782 19610
rect 13834 19558 13846 19610
rect 13898 19558 13910 19610
rect 13962 19558 13974 19610
rect 14026 19558 16782 19610
rect 16834 19558 16846 19610
rect 16898 19558 16910 19610
rect 16962 19558 16974 19610
rect 17026 19558 19782 19610
rect 19834 19558 19846 19610
rect 19898 19558 19910 19610
rect 19962 19558 19974 19610
rect 20026 19558 22782 19610
rect 22834 19558 22846 19610
rect 22898 19558 22910 19610
rect 22962 19558 22974 19610
rect 23026 19558 25782 19610
rect 25834 19558 25846 19610
rect 25898 19558 25910 19610
rect 25962 19558 25974 19610
rect 26026 19558 28336 19610
rect 1104 19536 28336 19558
rect 1104 19066 28336 19088
rect 1104 19014 3282 19066
rect 3334 19014 3346 19066
rect 3398 19014 3410 19066
rect 3462 19014 3474 19066
rect 3526 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 6410 19066
rect 6462 19014 6474 19066
rect 6526 19014 9282 19066
rect 9334 19014 9346 19066
rect 9398 19014 9410 19066
rect 9462 19014 9474 19066
rect 9526 19014 12282 19066
rect 12334 19014 12346 19066
rect 12398 19014 12410 19066
rect 12462 19014 12474 19066
rect 12526 19014 15282 19066
rect 15334 19014 15346 19066
rect 15398 19014 15410 19066
rect 15462 19014 15474 19066
rect 15526 19014 18282 19066
rect 18334 19014 18346 19066
rect 18398 19014 18410 19066
rect 18462 19014 18474 19066
rect 18526 19014 21282 19066
rect 21334 19014 21346 19066
rect 21398 19014 21410 19066
rect 21462 19014 21474 19066
rect 21526 19014 24282 19066
rect 24334 19014 24346 19066
rect 24398 19014 24410 19066
rect 24462 19014 24474 19066
rect 24526 19014 27282 19066
rect 27334 19014 27346 19066
rect 27398 19014 27410 19066
rect 27462 19014 27474 19066
rect 27526 19014 28336 19066
rect 1104 18992 28336 19014
rect 1104 18522 28336 18544
rect 1104 18470 1782 18522
rect 1834 18470 1846 18522
rect 1898 18470 1910 18522
rect 1962 18470 1974 18522
rect 2026 18470 4782 18522
rect 4834 18470 4846 18522
rect 4898 18470 4910 18522
rect 4962 18470 4974 18522
rect 5026 18470 7782 18522
rect 7834 18470 7846 18522
rect 7898 18470 7910 18522
rect 7962 18470 7974 18522
rect 8026 18470 10782 18522
rect 10834 18470 10846 18522
rect 10898 18470 10910 18522
rect 10962 18470 10974 18522
rect 11026 18470 13782 18522
rect 13834 18470 13846 18522
rect 13898 18470 13910 18522
rect 13962 18470 13974 18522
rect 14026 18470 16782 18522
rect 16834 18470 16846 18522
rect 16898 18470 16910 18522
rect 16962 18470 16974 18522
rect 17026 18470 19782 18522
rect 19834 18470 19846 18522
rect 19898 18470 19910 18522
rect 19962 18470 19974 18522
rect 20026 18470 22782 18522
rect 22834 18470 22846 18522
rect 22898 18470 22910 18522
rect 22962 18470 22974 18522
rect 23026 18470 25782 18522
rect 25834 18470 25846 18522
rect 25898 18470 25910 18522
rect 25962 18470 25974 18522
rect 26026 18470 28336 18522
rect 1104 18448 28336 18470
rect 1104 17978 28336 18000
rect 1104 17926 3282 17978
rect 3334 17926 3346 17978
rect 3398 17926 3410 17978
rect 3462 17926 3474 17978
rect 3526 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 6410 17978
rect 6462 17926 6474 17978
rect 6526 17926 9282 17978
rect 9334 17926 9346 17978
rect 9398 17926 9410 17978
rect 9462 17926 9474 17978
rect 9526 17926 12282 17978
rect 12334 17926 12346 17978
rect 12398 17926 12410 17978
rect 12462 17926 12474 17978
rect 12526 17926 15282 17978
rect 15334 17926 15346 17978
rect 15398 17926 15410 17978
rect 15462 17926 15474 17978
rect 15526 17926 18282 17978
rect 18334 17926 18346 17978
rect 18398 17926 18410 17978
rect 18462 17926 18474 17978
rect 18526 17926 21282 17978
rect 21334 17926 21346 17978
rect 21398 17926 21410 17978
rect 21462 17926 21474 17978
rect 21526 17926 24282 17978
rect 24334 17926 24346 17978
rect 24398 17926 24410 17978
rect 24462 17926 24474 17978
rect 24526 17926 27282 17978
rect 27334 17926 27346 17978
rect 27398 17926 27410 17978
rect 27462 17926 27474 17978
rect 27526 17926 28336 17978
rect 1104 17904 28336 17926
rect 1104 17434 28336 17456
rect 1104 17382 1782 17434
rect 1834 17382 1846 17434
rect 1898 17382 1910 17434
rect 1962 17382 1974 17434
rect 2026 17382 4782 17434
rect 4834 17382 4846 17434
rect 4898 17382 4910 17434
rect 4962 17382 4974 17434
rect 5026 17382 7782 17434
rect 7834 17382 7846 17434
rect 7898 17382 7910 17434
rect 7962 17382 7974 17434
rect 8026 17382 10782 17434
rect 10834 17382 10846 17434
rect 10898 17382 10910 17434
rect 10962 17382 10974 17434
rect 11026 17382 13782 17434
rect 13834 17382 13846 17434
rect 13898 17382 13910 17434
rect 13962 17382 13974 17434
rect 14026 17382 16782 17434
rect 16834 17382 16846 17434
rect 16898 17382 16910 17434
rect 16962 17382 16974 17434
rect 17026 17382 19782 17434
rect 19834 17382 19846 17434
rect 19898 17382 19910 17434
rect 19962 17382 19974 17434
rect 20026 17382 22782 17434
rect 22834 17382 22846 17434
rect 22898 17382 22910 17434
rect 22962 17382 22974 17434
rect 23026 17382 25782 17434
rect 25834 17382 25846 17434
rect 25898 17382 25910 17434
rect 25962 17382 25974 17434
rect 26026 17382 28336 17434
rect 1104 17360 28336 17382
rect 1104 16890 28336 16912
rect 1104 16838 3282 16890
rect 3334 16838 3346 16890
rect 3398 16838 3410 16890
rect 3462 16838 3474 16890
rect 3526 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 6410 16890
rect 6462 16838 6474 16890
rect 6526 16838 9282 16890
rect 9334 16838 9346 16890
rect 9398 16838 9410 16890
rect 9462 16838 9474 16890
rect 9526 16838 12282 16890
rect 12334 16838 12346 16890
rect 12398 16838 12410 16890
rect 12462 16838 12474 16890
rect 12526 16838 15282 16890
rect 15334 16838 15346 16890
rect 15398 16838 15410 16890
rect 15462 16838 15474 16890
rect 15526 16838 18282 16890
rect 18334 16838 18346 16890
rect 18398 16838 18410 16890
rect 18462 16838 18474 16890
rect 18526 16838 21282 16890
rect 21334 16838 21346 16890
rect 21398 16838 21410 16890
rect 21462 16838 21474 16890
rect 21526 16838 24282 16890
rect 24334 16838 24346 16890
rect 24398 16838 24410 16890
rect 24462 16838 24474 16890
rect 24526 16838 27282 16890
rect 27334 16838 27346 16890
rect 27398 16838 27410 16890
rect 27462 16838 27474 16890
rect 27526 16838 28336 16890
rect 1104 16816 28336 16838
rect 14734 16668 14740 16720
rect 14792 16708 14798 16720
rect 16761 16711 16819 16717
rect 16761 16708 16773 16711
rect 14792 16680 16773 16708
rect 14792 16668 14798 16680
rect 16761 16677 16773 16680
rect 16807 16677 16819 16711
rect 16761 16671 16819 16677
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16572 14243 16575
rect 14274 16572 14280 16584
rect 14231 16544 14280 16572
rect 14231 16541 14243 16544
rect 14185 16535 14243 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 16298 16572 16304 16584
rect 16163 16544 16304 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16298 16532 16304 16544
rect 16356 16532 16362 16584
rect 16482 16572 16488 16584
rect 16443 16544 16488 16572
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17126 16572 17132 16584
rect 16899 16544 17132 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 14366 16436 14372 16448
rect 14327 16408 14372 16436
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 15565 16439 15623 16445
rect 15565 16405 15577 16439
rect 15611 16436 15623 16439
rect 16114 16436 16120 16448
rect 15611 16408 16120 16436
rect 15611 16405 15623 16408
rect 15565 16399 15623 16405
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 1104 16346 28336 16368
rect 1104 16294 1782 16346
rect 1834 16294 1846 16346
rect 1898 16294 1910 16346
rect 1962 16294 1974 16346
rect 2026 16294 4782 16346
rect 4834 16294 4846 16346
rect 4898 16294 4910 16346
rect 4962 16294 4974 16346
rect 5026 16294 7782 16346
rect 7834 16294 7846 16346
rect 7898 16294 7910 16346
rect 7962 16294 7974 16346
rect 8026 16294 10782 16346
rect 10834 16294 10846 16346
rect 10898 16294 10910 16346
rect 10962 16294 10974 16346
rect 11026 16294 13782 16346
rect 13834 16294 13846 16346
rect 13898 16294 13910 16346
rect 13962 16294 13974 16346
rect 14026 16294 16782 16346
rect 16834 16294 16846 16346
rect 16898 16294 16910 16346
rect 16962 16294 16974 16346
rect 17026 16294 19782 16346
rect 19834 16294 19846 16346
rect 19898 16294 19910 16346
rect 19962 16294 19974 16346
rect 20026 16294 22782 16346
rect 22834 16294 22846 16346
rect 22898 16294 22910 16346
rect 22962 16294 22974 16346
rect 23026 16294 25782 16346
rect 25834 16294 25846 16346
rect 25898 16294 25910 16346
rect 25962 16294 25974 16346
rect 26026 16294 28336 16346
rect 1104 16272 28336 16294
rect 14185 16235 14243 16241
rect 14185 16201 14197 16235
rect 14231 16232 14243 16235
rect 14366 16232 14372 16244
rect 14231 16204 14372 16232
rect 14231 16201 14243 16204
rect 14185 16195 14243 16201
rect 14366 16192 14372 16204
rect 14424 16232 14430 16244
rect 14424 16204 15240 16232
rect 14424 16192 14430 16204
rect 14642 16164 14648 16176
rect 14476 16136 14648 16164
rect 14476 16105 14504 16136
rect 14642 16124 14648 16136
rect 14700 16124 14706 16176
rect 14734 16124 14740 16176
rect 14792 16164 14798 16176
rect 14792 16136 14837 16164
rect 15212 16136 15240 16204
rect 16298 16192 16304 16244
rect 16356 16232 16362 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16356 16204 16773 16232
rect 16356 16192 16362 16204
rect 16761 16201 16773 16204
rect 16807 16232 16819 16235
rect 17954 16232 17960 16244
rect 16807 16204 17960 16232
rect 16807 16201 16819 16204
rect 16761 16195 16819 16201
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 14792 16124 14798 16136
rect 14461 16099 14519 16105
rect 14461 16065 14473 16099
rect 14507 16065 14519 16099
rect 19886 16096 19892 16108
rect 19847 16068 19892 16096
rect 14461 16059 14519 16065
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 16114 15988 16120 16040
rect 16172 16028 16178 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 16172 16000 16497 16028
rect 16172 15988 16178 16000
rect 16485 15997 16497 16000
rect 16531 15997 16543 16031
rect 16485 15991 16543 15997
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 19245 16031 19303 16037
rect 19245 16028 19257 16031
rect 18196 16000 19257 16028
rect 18196 15988 18202 16000
rect 19245 15997 19257 16000
rect 19291 16028 19303 16031
rect 19610 16028 19616 16040
rect 19291 16000 19616 16028
rect 19291 15997 19303 16000
rect 19245 15991 19303 15997
rect 19610 15988 19616 16000
rect 19668 15988 19674 16040
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 17126 15892 17132 15904
rect 13872 15864 13917 15892
rect 17087 15864 17132 15892
rect 13872 15852 13878 15864
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 1104 15802 28336 15824
rect 1104 15750 3282 15802
rect 3334 15750 3346 15802
rect 3398 15750 3410 15802
rect 3462 15750 3474 15802
rect 3526 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 6410 15802
rect 6462 15750 6474 15802
rect 6526 15750 9282 15802
rect 9334 15750 9346 15802
rect 9398 15750 9410 15802
rect 9462 15750 9474 15802
rect 9526 15750 12282 15802
rect 12334 15750 12346 15802
rect 12398 15750 12410 15802
rect 12462 15750 12474 15802
rect 12526 15750 15282 15802
rect 15334 15750 15346 15802
rect 15398 15750 15410 15802
rect 15462 15750 15474 15802
rect 15526 15750 18282 15802
rect 18334 15750 18346 15802
rect 18398 15750 18410 15802
rect 18462 15750 18474 15802
rect 18526 15750 21282 15802
rect 21334 15750 21346 15802
rect 21398 15750 21410 15802
rect 21462 15750 21474 15802
rect 21526 15750 24282 15802
rect 24334 15750 24346 15802
rect 24398 15750 24410 15802
rect 24462 15750 24474 15802
rect 24526 15750 27282 15802
rect 27334 15750 27346 15802
rect 27398 15750 27410 15802
rect 27462 15750 27474 15802
rect 27526 15750 28336 15802
rect 1104 15728 28336 15750
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 16482 15648 16488 15660
rect 16540 15688 16546 15700
rect 17405 15691 17463 15697
rect 17405 15688 17417 15691
rect 16540 15660 17417 15688
rect 16540 15648 16546 15660
rect 17405 15657 17417 15660
rect 17451 15657 17463 15691
rect 17405 15651 17463 15657
rect 13814 15552 13820 15564
rect 13786 15512 13820 15552
rect 13872 15552 13878 15564
rect 14274 15552 14280 15564
rect 13872 15524 14280 15552
rect 13872 15512 13878 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 14369 15555 14427 15561
rect 14369 15521 14381 15555
rect 14415 15552 14427 15555
rect 17126 15552 17132 15564
rect 14415 15524 17132 15552
rect 14415 15521 14427 15524
rect 14369 15515 14427 15521
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 17460 15524 18061 15552
rect 17460 15512 17466 15524
rect 18049 15521 18061 15524
rect 18095 15521 18107 15555
rect 18049 15515 18107 15521
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19705 15555 19763 15561
rect 19705 15552 19717 15555
rect 19484 15524 19717 15552
rect 19484 15512 19490 15524
rect 19705 15521 19717 15524
rect 19751 15552 19763 15555
rect 19886 15552 19892 15564
rect 19751 15524 19892 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 19886 15512 19892 15524
rect 19944 15552 19950 15564
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 19944 15524 20085 15552
rect 19944 15512 19950 15524
rect 20073 15521 20085 15524
rect 20119 15552 20131 15555
rect 20714 15552 20720 15564
rect 20119 15524 20720 15552
rect 20119 15521 20131 15524
rect 20073 15515 20131 15521
rect 20714 15512 20720 15524
rect 20772 15552 20778 15564
rect 23109 15555 23167 15561
rect 23109 15552 23121 15555
rect 20772 15524 23121 15552
rect 20772 15512 20778 15524
rect 23109 15521 23121 15524
rect 23155 15521 23167 15555
rect 23109 15515 23167 15521
rect 12802 15484 12808 15496
rect 12763 15456 12808 15484
rect 12802 15444 12808 15456
rect 12860 15484 12866 15496
rect 13786 15484 13814 15512
rect 12860 15456 13814 15484
rect 14001 15487 14059 15493
rect 12860 15444 12866 15456
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 14550 15484 14556 15496
rect 14047 15456 14556 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 16114 15484 16120 15496
rect 16075 15456 16120 15484
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17586 15484 17592 15496
rect 17547 15456 17592 15484
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17736 15456 17785 15484
rect 17736 15444 17742 15456
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 18138 15484 18144 15496
rect 18099 15456 18144 15484
rect 17773 15447 17831 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 19150 15484 19156 15496
rect 19111 15456 19156 15484
rect 19150 15444 19156 15456
rect 19208 15444 19214 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 13541 15419 13599 15425
rect 13541 15385 13553 15419
rect 13587 15416 13599 15419
rect 13817 15419 13875 15425
rect 13817 15416 13829 15419
rect 13587 15388 13829 15416
rect 13587 15385 13599 15388
rect 13541 15379 13599 15385
rect 13817 15385 13829 15388
rect 13863 15416 13875 15419
rect 13863 15388 15976 15416
rect 13863 15385 13875 15388
rect 13817 15379 13875 15385
rect 15948 15360 15976 15388
rect 21266 15376 21272 15428
rect 21324 15416 21330 15428
rect 21361 15419 21419 15425
rect 21361 15416 21373 15419
rect 21324 15388 21373 15416
rect 21324 15376 21330 15388
rect 21361 15385 21373 15388
rect 21407 15385 21419 15419
rect 21361 15379 21419 15385
rect 21910 15376 21916 15428
rect 21968 15376 21974 15428
rect 12986 15348 12992 15360
rect 12947 15320 12992 15348
rect 12986 15308 12992 15320
rect 13044 15348 13050 15360
rect 13354 15348 13360 15360
rect 13044 15320 13360 15348
rect 13044 15308 13050 15320
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 14642 15348 14648 15360
rect 14603 15320 14648 15348
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 15930 15348 15936 15360
rect 15891 15320 15936 15348
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 19337 15351 19395 15357
rect 19337 15317 19349 15351
rect 19383 15348 19395 15351
rect 19518 15348 19524 15360
rect 19383 15320 19524 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 1104 15258 28336 15280
rect 1104 15206 1782 15258
rect 1834 15206 1846 15258
rect 1898 15206 1910 15258
rect 1962 15206 1974 15258
rect 2026 15206 4782 15258
rect 4834 15206 4846 15258
rect 4898 15206 4910 15258
rect 4962 15206 4974 15258
rect 5026 15206 7782 15258
rect 7834 15206 7846 15258
rect 7898 15206 7910 15258
rect 7962 15206 7974 15258
rect 8026 15206 10782 15258
rect 10834 15206 10846 15258
rect 10898 15206 10910 15258
rect 10962 15206 10974 15258
rect 11026 15206 13782 15258
rect 13834 15206 13846 15258
rect 13898 15206 13910 15258
rect 13962 15206 13974 15258
rect 14026 15206 16782 15258
rect 16834 15206 16846 15258
rect 16898 15206 16910 15258
rect 16962 15206 16974 15258
rect 17026 15206 19782 15258
rect 19834 15206 19846 15258
rect 19898 15206 19910 15258
rect 19962 15206 19974 15258
rect 20026 15206 22782 15258
rect 22834 15206 22846 15258
rect 22898 15206 22910 15258
rect 22962 15206 22974 15258
rect 23026 15206 25782 15258
rect 25834 15206 25846 15258
rect 25898 15206 25910 15258
rect 25962 15206 25974 15258
rect 26026 15206 28336 15258
rect 1104 15184 28336 15206
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15144 12127 15147
rect 12802 15144 12808 15156
rect 12115 15116 12808 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 14642 15144 14648 15156
rect 12912 15116 14648 15144
rect 12912 15076 12940 15116
rect 14642 15104 14648 15116
rect 14700 15104 14706 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14792 15116 14933 15144
rect 14792 15104 14798 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21082 15144 21088 15156
rect 21039 15116 21088 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 21637 15147 21695 15153
rect 21637 15113 21649 15147
rect 21683 15144 21695 15147
rect 21910 15144 21916 15156
rect 21683 15116 21916 15144
rect 21683 15113 21695 15116
rect 21637 15107 21695 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 12636 15048 12940 15076
rect 12636 14952 12664 15048
rect 13354 15036 13360 15088
rect 13412 15036 13418 15088
rect 17589 15079 17647 15085
rect 17589 15045 17601 15079
rect 17635 15076 17647 15079
rect 18138 15076 18144 15088
rect 17635 15048 18144 15076
rect 17635 15045 17647 15048
rect 17589 15039 17647 15045
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 18509 15079 18567 15085
rect 18509 15045 18521 15079
rect 18555 15076 18567 15079
rect 19150 15076 19156 15088
rect 18555 15048 19156 15076
rect 18555 15045 18567 15048
rect 18509 15039 18567 15045
rect 19150 15036 19156 15048
rect 19208 15076 19214 15088
rect 20346 15076 20352 15088
rect 19208 15048 20352 15076
rect 19208 15036 19214 15048
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 14240 14980 14657 15008
rect 14240 14968 14246 14980
rect 14645 14977 14657 14980
rect 14691 15008 14703 15011
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 14691 14980 15485 15008
rect 14691 14977 14703 14980
rect 14645 14971 14703 14977
rect 15473 14977 15485 14980
rect 15519 15008 15531 15011
rect 15746 15008 15752 15020
rect 15519 14980 15752 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 19426 15008 19432 15020
rect 19387 14980 19432 15008
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 19536 14980 19993 15008
rect 12618 14940 12624 14952
rect 12579 14912 12624 14940
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 12894 14940 12900 14952
rect 12855 14912 12900 14940
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 16485 14943 16543 14949
rect 16485 14909 16497 14943
rect 16531 14940 16543 14943
rect 17678 14940 17684 14952
rect 16531 14912 17684 14940
rect 16531 14909 16543 14912
rect 16485 14903 16543 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 18012 14912 19257 14940
rect 18012 14900 18018 14912
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 16853 14875 16911 14881
rect 16853 14841 16865 14875
rect 16899 14872 16911 14875
rect 17586 14872 17592 14884
rect 16899 14844 17592 14872
rect 16899 14841 16911 14844
rect 16853 14835 16911 14841
rect 17586 14832 17592 14844
rect 17644 14832 17650 14884
rect 18966 14832 18972 14884
rect 19024 14872 19030 14884
rect 19536 14872 19564 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 20162 15008 20168 15020
rect 20123 14980 20168 15008
rect 19981 14971 20039 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 15008 21511 15011
rect 21634 15008 21640 15020
rect 21499 14980 21640 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14940 20591 14943
rect 21174 14940 21180 14952
rect 20579 14912 21180 14940
rect 20579 14909 20591 14912
rect 20533 14903 20591 14909
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 19024 14844 19564 14872
rect 19024 14832 19030 14844
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 17221 14807 17279 14813
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 17402 14804 17408 14816
rect 17267 14776 17408 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 18874 14804 18880 14816
rect 18835 14776 18880 14804
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 1104 14714 28336 14736
rect 1104 14662 3282 14714
rect 3334 14662 3346 14714
rect 3398 14662 3410 14714
rect 3462 14662 3474 14714
rect 3526 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 6410 14714
rect 6462 14662 6474 14714
rect 6526 14662 9282 14714
rect 9334 14662 9346 14714
rect 9398 14662 9410 14714
rect 9462 14662 9474 14714
rect 9526 14662 12282 14714
rect 12334 14662 12346 14714
rect 12398 14662 12410 14714
rect 12462 14662 12474 14714
rect 12526 14662 15282 14714
rect 15334 14662 15346 14714
rect 15398 14662 15410 14714
rect 15462 14662 15474 14714
rect 15526 14662 18282 14714
rect 18334 14662 18346 14714
rect 18398 14662 18410 14714
rect 18462 14662 18474 14714
rect 18526 14662 21282 14714
rect 21334 14662 21346 14714
rect 21398 14662 21410 14714
rect 21462 14662 21474 14714
rect 21526 14662 24282 14714
rect 24334 14662 24346 14714
rect 24398 14662 24410 14714
rect 24462 14662 24474 14714
rect 24526 14662 27282 14714
rect 27334 14662 27346 14714
rect 27398 14662 27410 14714
rect 27462 14662 27474 14714
rect 27526 14662 28336 14714
rect 1104 14640 28336 14662
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 14550 14600 14556 14612
rect 14148 14572 14556 14600
rect 14148 14560 14154 14572
rect 14550 14560 14556 14572
rect 14608 14600 14614 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14608 14572 14657 14600
rect 14608 14560 14614 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 17405 14603 17463 14609
rect 17405 14569 17417 14603
rect 17451 14600 17463 14603
rect 17586 14600 17592 14612
rect 17451 14572 17592 14600
rect 17451 14569 17463 14572
rect 17405 14563 17463 14569
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 18012 14572 18429 14600
rect 18012 14560 18018 14572
rect 18417 14569 18429 14572
rect 18463 14600 18475 14603
rect 20162 14600 20168 14612
rect 18463 14572 20168 14600
rect 18463 14569 18475 14572
rect 18417 14563 18475 14569
rect 20162 14560 20168 14572
rect 20220 14600 20226 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 20220 14572 20269 14600
rect 20220 14560 20226 14572
rect 20257 14569 20269 14572
rect 20303 14569 20315 14603
rect 21174 14600 21180 14612
rect 21135 14572 21180 14600
rect 20257 14563 20315 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 21545 14603 21603 14609
rect 21545 14569 21557 14603
rect 21591 14600 21603 14603
rect 21634 14600 21640 14612
rect 21591 14572 21640 14600
rect 21591 14569 21603 14572
rect 21545 14563 21603 14569
rect 21634 14560 21640 14572
rect 21692 14560 21698 14612
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14464 12311 14467
rect 12894 14464 12900 14476
rect 12299 14436 12900 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 14182 14464 14188 14476
rect 13004 14436 14188 14464
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11572 14368 11897 14396
rect 11572 14356 11578 14368
rect 11885 14365 11897 14368
rect 11931 14396 11943 14399
rect 13004 14396 13032 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14366 14424 14372 14476
rect 14424 14464 14430 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 14424 14436 15577 14464
rect 14424 14424 14430 14436
rect 15565 14433 15577 14436
rect 15611 14464 15623 14467
rect 15654 14464 15660 14476
rect 15611 14436 15660 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 15654 14424 15660 14436
rect 15712 14464 15718 14476
rect 16485 14467 16543 14473
rect 16485 14464 16497 14467
rect 15712 14436 16497 14464
rect 15712 14424 15718 14436
rect 16485 14433 16497 14436
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 19245 14467 19303 14473
rect 19245 14433 19257 14467
rect 19291 14464 19303 14467
rect 20254 14464 20260 14476
rect 19291 14436 20260 14464
rect 19291 14433 19303 14436
rect 19245 14427 19303 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 21082 14424 21088 14476
rect 21140 14464 21146 14476
rect 21910 14464 21916 14476
rect 21140 14436 21916 14464
rect 21140 14424 21146 14436
rect 21910 14424 21916 14436
rect 21968 14464 21974 14476
rect 22373 14467 22431 14473
rect 22373 14464 22385 14467
rect 21968 14436 22385 14464
rect 21968 14424 21974 14436
rect 22373 14433 22385 14436
rect 22419 14433 22431 14467
rect 22373 14427 22431 14433
rect 23842 14424 23848 14476
rect 23900 14464 23906 14476
rect 24397 14467 24455 14473
rect 24397 14464 24409 14467
rect 23900 14436 24409 14464
rect 23900 14424 23906 14436
rect 24397 14433 24409 14436
rect 24443 14433 24455 14467
rect 24397 14427 24455 14433
rect 13354 14396 13360 14408
rect 11931 14368 13032 14396
rect 13315 14368 13360 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 13538 14396 13544 14408
rect 13499 14368 13544 14396
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13688 14368 13737 14396
rect 13688 14356 13694 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 14277 14359 14335 14365
rect 12710 14288 12716 14340
rect 12768 14328 12774 14340
rect 14292 14328 14320 14359
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 15930 14396 15936 14408
rect 15795 14368 15936 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 15930 14356 15936 14368
rect 15988 14396 15994 14408
rect 16666 14396 16672 14408
rect 15988 14368 16672 14396
rect 15988 14356 15994 14368
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17586 14396 17592 14408
rect 17547 14368 17592 14396
rect 17586 14356 17592 14368
rect 17644 14356 17650 14408
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14396 18199 14399
rect 18966 14396 18972 14408
rect 18187 14368 18972 14396
rect 18187 14365 18199 14368
rect 18141 14359 18199 14365
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19668 14368 19809 14396
rect 19668 14356 19674 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20162 14396 20168 14408
rect 20027 14368 20168 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 12768 14300 14320 14328
rect 12768 14288 12774 14300
rect 11422 14220 11428 14272
rect 11480 14260 11486 14272
rect 12529 14263 12587 14269
rect 12529 14260 12541 14263
rect 11480 14232 12541 14260
rect 11480 14220 11486 14232
rect 12529 14229 12541 14232
rect 12575 14260 12587 14263
rect 12618 14260 12624 14272
rect 12575 14232 12624 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 14292 14260 14320 14300
rect 16209 14331 16267 14337
rect 16209 14297 16221 14331
rect 16255 14328 16267 14331
rect 16390 14328 16396 14340
rect 16255 14300 16396 14328
rect 16255 14297 16267 14300
rect 16209 14291 16267 14297
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 19812 14328 19840 14359
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20530 14328 20536 14340
rect 19812 14300 20536 14328
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 22646 14328 22652 14340
rect 22607 14300 22652 14328
rect 22646 14288 22652 14300
rect 22704 14288 22710 14340
rect 23106 14288 23112 14340
rect 23164 14288 23170 14340
rect 17770 14260 17776 14272
rect 14292 14232 17776 14260
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 19058 14260 19064 14272
rect 18971 14232 19064 14260
rect 19058 14220 19064 14232
rect 19116 14260 19122 14272
rect 19610 14260 19616 14272
rect 19116 14232 19616 14260
rect 19116 14220 19122 14232
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 1104 14170 28336 14192
rect 1104 14118 1782 14170
rect 1834 14118 1846 14170
rect 1898 14118 1910 14170
rect 1962 14118 1974 14170
rect 2026 14118 4782 14170
rect 4834 14118 4846 14170
rect 4898 14118 4910 14170
rect 4962 14118 4974 14170
rect 5026 14118 7782 14170
rect 7834 14118 7846 14170
rect 7898 14118 7910 14170
rect 7962 14118 7974 14170
rect 8026 14118 10782 14170
rect 10834 14118 10846 14170
rect 10898 14118 10910 14170
rect 10962 14118 10974 14170
rect 11026 14118 13782 14170
rect 13834 14118 13846 14170
rect 13898 14118 13910 14170
rect 13962 14118 13974 14170
rect 14026 14118 16782 14170
rect 16834 14118 16846 14170
rect 16898 14118 16910 14170
rect 16962 14118 16974 14170
rect 17026 14118 19782 14170
rect 19834 14118 19846 14170
rect 19898 14118 19910 14170
rect 19962 14118 19974 14170
rect 20026 14118 22782 14170
rect 22834 14118 22846 14170
rect 22898 14118 22910 14170
rect 22962 14118 22974 14170
rect 23026 14118 25782 14170
rect 25834 14118 25846 14170
rect 25898 14118 25910 14170
rect 25962 14118 25974 14170
rect 26026 14118 28336 14170
rect 1104 14096 28336 14118
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 12986 14056 12992 14068
rect 12759 14028 12992 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13081 14059 13139 14065
rect 13081 14025 13093 14059
rect 13127 14056 13139 14059
rect 13262 14056 13268 14068
rect 13127 14028 13268 14056
rect 13127 14025 13139 14028
rect 13081 14019 13139 14025
rect 13262 14016 13268 14028
rect 13320 14056 13326 14068
rect 13630 14056 13636 14068
rect 13320 14028 13636 14056
rect 13320 14016 13326 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15470 14056 15476 14068
rect 15151 14028 15476 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 15470 14016 15476 14028
rect 15528 14056 15534 14068
rect 17310 14056 17316 14068
rect 15528 14028 17316 14056
rect 15528 14016 15534 14028
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18966 14056 18972 14068
rect 18927 14028 18972 14056
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19150 14056 19156 14068
rect 19076 14028 19156 14056
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13988 12127 13991
rect 13354 13988 13360 14000
rect 12115 13960 13360 13988
rect 12115 13957 12127 13960
rect 12069 13951 12127 13957
rect 13354 13948 13360 13960
rect 13412 13988 13418 14000
rect 13541 13991 13599 13997
rect 13541 13988 13553 13991
rect 13412 13960 13553 13988
rect 13412 13948 13418 13960
rect 13541 13957 13553 13960
rect 13587 13957 13599 13991
rect 15562 13988 15568 14000
rect 13541 13951 13599 13957
rect 14476 13960 15568 13988
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 8757 13923 8815 13929
rect 8757 13920 8769 13923
rect 8536 13892 8769 13920
rect 8536 13880 8542 13892
rect 8757 13889 8769 13892
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13504 13892 14013 13920
rect 13504 13880 13510 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14366 13920 14372 13932
rect 14327 13892 14372 13920
rect 14001 13883 14059 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 14476 13929 14504 13960
rect 15562 13948 15568 13960
rect 15620 13988 15626 14000
rect 17037 13991 17095 13997
rect 15620 13960 16252 13988
rect 15620 13948 15626 13960
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14461 13883 14519 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 15746 13920 15752 13932
rect 15703 13892 15752 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 16224 13920 16252 13960
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 17586 13988 17592 14000
rect 17083 13960 17592 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 17681 13991 17739 13997
rect 17681 13957 17693 13991
rect 17727 13988 17739 13991
rect 19076 13988 19104 14028
rect 19150 14016 19156 14028
rect 19208 14056 19214 14068
rect 19208 14028 19334 14056
rect 19208 14016 19214 14028
rect 17727 13960 19104 13988
rect 19306 13988 19334 14028
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 19484 14028 20177 14056
rect 19484 14016 19490 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 19306 13960 19748 13988
rect 17727 13957 17739 13960
rect 17681 13951 17739 13957
rect 17696 13920 17724 13951
rect 16224 13892 17724 13920
rect 18874 13880 18880 13932
rect 18932 13920 18938 13932
rect 19720 13929 19748 13960
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 18932 13892 19349 13920
rect 18932 13880 18938 13892
rect 19337 13889 19349 13892
rect 19383 13889 19395 13923
rect 19337 13883 19395 13889
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13889 19763 13923
rect 20180 13920 20208 14019
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 20404 14028 21465 14056
rect 20404 14016 20410 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 23106 14056 23112 14068
rect 23067 14028 23112 14056
rect 21453 14019 21511 14025
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 20254 13948 20260 14000
rect 20312 13988 20318 14000
rect 20312 13960 21312 13988
rect 20312 13948 20318 13960
rect 20990 13920 20996 13932
rect 20180 13892 20996 13920
rect 19705 13883 19763 13889
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 15381 13855 15439 13861
rect 15381 13852 15393 13855
rect 13596 13824 15393 13852
rect 13596 13812 13602 13824
rect 15381 13821 15393 13824
rect 15427 13852 15439 13855
rect 16114 13852 16120 13864
rect 15427 13824 16120 13852
rect 15427 13821 15439 13824
rect 15381 13815 15439 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 16666 13852 16672 13864
rect 16531 13824 16672 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 19153 13855 19211 13861
rect 19153 13852 19165 13855
rect 17460 13824 19165 13852
rect 17460 13812 17466 13824
rect 19153 13821 19165 13824
rect 19199 13821 19211 13855
rect 19153 13815 19211 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19426 13852 19432 13864
rect 19291 13824 19432 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19610 13852 19616 13864
rect 19571 13824 19616 13852
rect 19610 13812 19616 13824
rect 19668 13812 19674 13864
rect 20070 13744 20076 13796
rect 20128 13784 20134 13796
rect 20272 13784 20300 13892
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 21284 13929 21312 13960
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 20530 13852 20536 13864
rect 20491 13824 20536 13852
rect 20530 13812 20536 13824
rect 20588 13852 20594 13864
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20588 13824 21097 13852
rect 20588 13812 20594 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 20128 13756 20300 13784
rect 20128 13744 20134 13756
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22373 13787 22431 13793
rect 22373 13784 22385 13787
rect 22152 13756 22385 13784
rect 22152 13744 22158 13756
rect 22373 13753 22385 13756
rect 22419 13753 22431 13787
rect 22373 13747 22431 13753
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8904 13688 8953 13716
rect 8904 13676 8910 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 8941 13679 8999 13685
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 11514 13716 11520 13728
rect 11379 13688 11520 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11698 13716 11704 13728
rect 11659 13688 11704 13716
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 15838 13716 15844 13728
rect 15799 13688 15844 13716
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 18417 13719 18475 13725
rect 18417 13685 18429 13719
rect 18463 13716 18475 13719
rect 18690 13716 18696 13728
rect 18463 13688 18696 13716
rect 18463 13685 18475 13688
rect 18417 13679 18475 13685
rect 18690 13676 18696 13688
rect 18748 13716 18754 13728
rect 20162 13716 20168 13728
rect 18748 13688 20168 13716
rect 18748 13676 18754 13688
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 22646 13676 22652 13728
rect 22704 13716 22710 13728
rect 22741 13719 22799 13725
rect 22741 13716 22753 13719
rect 22704 13688 22753 13716
rect 22704 13676 22710 13688
rect 22741 13685 22753 13688
rect 22787 13685 22799 13719
rect 22741 13679 22799 13685
rect 1104 13626 28336 13648
rect 1104 13574 3282 13626
rect 3334 13574 3346 13626
rect 3398 13574 3410 13626
rect 3462 13574 3474 13626
rect 3526 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 6410 13626
rect 6462 13574 6474 13626
rect 6526 13574 9282 13626
rect 9334 13574 9346 13626
rect 9398 13574 9410 13626
rect 9462 13574 9474 13626
rect 9526 13574 12282 13626
rect 12334 13574 12346 13626
rect 12398 13574 12410 13626
rect 12462 13574 12474 13626
rect 12526 13574 15282 13626
rect 15334 13574 15346 13626
rect 15398 13574 15410 13626
rect 15462 13574 15474 13626
rect 15526 13574 18282 13626
rect 18334 13574 18346 13626
rect 18398 13574 18410 13626
rect 18462 13574 18474 13626
rect 18526 13574 21282 13626
rect 21334 13574 21346 13626
rect 21398 13574 21410 13626
rect 21462 13574 21474 13626
rect 21526 13574 24282 13626
rect 24334 13574 24346 13626
rect 24398 13574 24410 13626
rect 24462 13574 24474 13626
rect 24526 13574 27282 13626
rect 27334 13574 27346 13626
rect 27398 13574 27410 13626
rect 27462 13574 27474 13626
rect 27526 13574 28336 13626
rect 1104 13552 28336 13574
rect 11514 13512 11520 13524
rect 11475 13484 11520 13512
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 12253 13515 12311 13521
rect 12253 13481 12265 13515
rect 12299 13512 12311 13515
rect 12710 13512 12716 13524
rect 12299 13484 12716 13512
rect 12299 13481 12311 13484
rect 12253 13475 12311 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 15746 13512 15752 13524
rect 15707 13484 15752 13512
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 18233 13515 18291 13521
rect 18233 13481 18245 13515
rect 18279 13512 18291 13515
rect 18874 13512 18880 13524
rect 18279 13484 18880 13512
rect 18279 13481 18291 13484
rect 18233 13475 18291 13481
rect 18874 13472 18880 13484
rect 18932 13512 18938 13524
rect 20073 13515 20131 13521
rect 20073 13512 20085 13515
rect 18932 13484 20085 13512
rect 18932 13472 18938 13484
rect 20073 13481 20085 13484
rect 20119 13512 20131 13515
rect 20254 13512 20260 13524
rect 20119 13484 20260 13512
rect 20119 13481 20131 13484
rect 20073 13475 20131 13481
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20530 13512 20536 13524
rect 20491 13484 20536 13512
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 20990 13472 20996 13524
rect 21048 13512 21054 13524
rect 21545 13515 21603 13521
rect 21545 13512 21557 13515
rect 21048 13484 21557 13512
rect 21048 13472 21054 13484
rect 21545 13481 21557 13484
rect 21591 13481 21603 13515
rect 21545 13475 21603 13481
rect 12621 13447 12679 13453
rect 12621 13413 12633 13447
rect 12667 13444 12679 13447
rect 14366 13444 14372 13456
rect 12667 13416 14372 13444
rect 12667 13413 12679 13416
rect 12621 13407 12679 13413
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 14737 13447 14795 13453
rect 14737 13413 14749 13447
rect 14783 13444 14795 13447
rect 15562 13444 15568 13456
rect 14783 13416 15568 13444
rect 14783 13413 14795 13416
rect 14737 13407 14795 13413
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 18969 13447 19027 13453
rect 18969 13413 18981 13447
rect 19015 13444 19027 13447
rect 19150 13444 19156 13456
rect 19015 13416 19156 13444
rect 19015 13413 19027 13416
rect 18969 13407 19027 13413
rect 19150 13404 19156 13416
rect 19208 13404 19214 13456
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19613 13447 19671 13453
rect 19613 13444 19625 13447
rect 19484 13416 19625 13444
rect 19484 13404 19490 13416
rect 19613 13413 19625 13416
rect 19659 13444 19671 13447
rect 21269 13447 21327 13453
rect 21269 13444 21281 13447
rect 19659 13416 21281 13444
rect 19659 13413 19671 13416
rect 19613 13407 19671 13413
rect 21269 13413 21281 13416
rect 21315 13413 21327 13447
rect 21269 13407 21327 13413
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13376 13047 13379
rect 13446 13376 13452 13388
rect 13035 13348 13452 13376
rect 13035 13345 13047 13348
rect 12989 13339 13047 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 13630 13336 13636 13388
rect 13688 13376 13694 13388
rect 13998 13376 14004 13388
rect 13688 13348 14004 13376
rect 13688 13336 13694 13348
rect 13998 13336 14004 13348
rect 14056 13336 14062 13388
rect 14182 13376 14188 13388
rect 14143 13348 14188 13376
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 16114 13376 16120 13388
rect 15887 13348 16120 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 17037 13379 17095 13385
rect 17037 13345 17049 13379
rect 17083 13376 17095 13379
rect 17218 13376 17224 13388
rect 17083 13348 17224 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 13817 13311 13875 13317
rect 13817 13277 13829 13311
rect 13863 13277 13875 13311
rect 14016 13308 14044 13336
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 14016 13280 14105 13308
rect 13817 13271 13875 13277
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 13832 13240 13860 13271
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 15620 13311 15678 13317
rect 15620 13308 15632 13311
rect 14608 13280 15632 13308
rect 14608 13268 14614 13280
rect 15620 13277 15632 13280
rect 15666 13277 15678 13311
rect 15620 13271 15678 13277
rect 17126 13268 17132 13320
rect 17184 13308 17190 13320
rect 19153 13311 19211 13317
rect 17184 13280 17229 13308
rect 17184 13268 17190 13280
rect 19153 13277 19165 13311
rect 19199 13308 19211 13311
rect 19518 13308 19524 13320
rect 19199 13280 19524 13308
rect 19199 13277 19211 13280
rect 19153 13271 19211 13277
rect 19518 13268 19524 13280
rect 19576 13268 19582 13320
rect 21082 13308 21088 13320
rect 21043 13280 21088 13308
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 14826 13240 14832 13252
rect 13832 13212 14832 13240
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 15473 13243 15531 13249
rect 15473 13240 15485 13243
rect 15160 13212 15485 13240
rect 15160 13200 15166 13212
rect 15473 13209 15485 13212
rect 15519 13209 15531 13243
rect 15473 13203 15531 13209
rect 16761 13243 16819 13249
rect 16761 13209 16773 13243
rect 16807 13240 16819 13243
rect 17144 13240 17172 13268
rect 17586 13240 17592 13252
rect 16807 13212 17172 13240
rect 17499 13212 17592 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 17586 13200 17592 13212
rect 17644 13240 17650 13252
rect 18782 13240 18788 13252
rect 17644 13212 18788 13240
rect 17644 13200 17650 13212
rect 18782 13200 18788 13212
rect 18840 13200 18846 13252
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 8478 13172 8484 13184
rect 8168 13144 8484 13172
rect 8168 13132 8174 13144
rect 8478 13132 8484 13144
rect 8536 13172 8542 13184
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8536 13144 8769 13172
rect 8536 13132 8542 13144
rect 8757 13141 8769 13144
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11756 13144 11897 13172
rect 11756 13132 11762 13144
rect 11885 13141 11897 13144
rect 11931 13172 11943 13175
rect 13538 13172 13544 13184
rect 11931 13144 13544 13172
rect 11931 13141 11943 13144
rect 11885 13135 11943 13141
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 16117 13175 16175 13181
rect 16117 13141 16129 13175
rect 16163 13172 16175 13175
rect 20990 13172 20996 13184
rect 16163 13144 20996 13172
rect 16163 13141 16175 13144
rect 16117 13135 16175 13141
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 23750 13172 23756 13184
rect 23711 13144 23756 13172
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 1104 13082 28336 13104
rect 1104 13030 1782 13082
rect 1834 13030 1846 13082
rect 1898 13030 1910 13082
rect 1962 13030 1974 13082
rect 2026 13030 4782 13082
rect 4834 13030 4846 13082
rect 4898 13030 4910 13082
rect 4962 13030 4974 13082
rect 5026 13030 7782 13082
rect 7834 13030 7846 13082
rect 7898 13030 7910 13082
rect 7962 13030 7974 13082
rect 8026 13030 10782 13082
rect 10834 13030 10846 13082
rect 10898 13030 10910 13082
rect 10962 13030 10974 13082
rect 11026 13030 13782 13082
rect 13834 13030 13846 13082
rect 13898 13030 13910 13082
rect 13962 13030 13974 13082
rect 14026 13030 16782 13082
rect 16834 13030 16846 13082
rect 16898 13030 16910 13082
rect 16962 13030 16974 13082
rect 17026 13030 19782 13082
rect 19834 13030 19846 13082
rect 19898 13030 19910 13082
rect 19962 13030 19974 13082
rect 20026 13030 22782 13082
rect 22834 13030 22846 13082
rect 22898 13030 22910 13082
rect 22962 13030 22974 13082
rect 23026 13030 25782 13082
rect 25834 13030 25846 13082
rect 25898 13030 25910 13082
rect 25962 13030 25974 13082
rect 26026 13030 28336 13082
rect 1104 13008 28336 13030
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11572 12940 11621 12968
rect 11572 12928 11578 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 11609 12931 11667 12937
rect 11624 12900 11652 12931
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 15473 12971 15531 12977
rect 13320 12940 13492 12968
rect 13320 12928 13326 12940
rect 11624 12872 13308 12900
rect 9122 12832 9128 12844
rect 9083 12804 9128 12832
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 13280 12841 13308 12872
rect 13464 12841 13492 12940
rect 15473 12937 15485 12971
rect 15519 12968 15531 12971
rect 15562 12968 15568 12980
rect 15519 12940 15568 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 18509 12971 18567 12977
rect 18509 12968 18521 12971
rect 17184 12940 18521 12968
rect 17184 12928 17190 12940
rect 18509 12937 18521 12940
rect 18555 12937 18567 12971
rect 19058 12968 19064 12980
rect 19019 12940 19064 12968
rect 18509 12931 18567 12937
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19518 12968 19524 12980
rect 19479 12940 19524 12968
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 17144 12900 17172 12928
rect 16592 12872 17172 12900
rect 18233 12903 18291 12909
rect 16592 12844 16620 12872
rect 18233 12869 18245 12903
rect 18279 12900 18291 12903
rect 18598 12900 18604 12912
rect 18279 12872 18604 12900
rect 18279 12869 18291 12872
rect 18233 12863 18291 12869
rect 18598 12860 18604 12872
rect 18656 12900 18662 12912
rect 19536 12900 19564 12928
rect 18656 12872 19564 12900
rect 18656 12860 18662 12872
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13265 12835 13323 12841
rect 13127 12804 13216 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 8662 12764 8668 12776
rect 8623 12736 8668 12764
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 11848 12736 12633 12764
rect 11848 12724 11854 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 13188 12696 13216 12804
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12801 13507 12835
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13449 12795 13507 12801
rect 13556 12804 14013 12832
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 13556 12764 13584 12804
rect 14001 12801 14013 12804
rect 14047 12832 14059 12835
rect 14182 12832 14188 12844
rect 14047 12804 14188 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 16574 12832 16580 12844
rect 16487 12804 16580 12832
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16816 12804 16865 12832
rect 16816 12792 16822 12804
rect 16853 12801 16865 12804
rect 16899 12832 16911 12835
rect 17402 12832 17408 12844
rect 16899 12804 17408 12832
rect 16899 12801 16911 12804
rect 16853 12795 16911 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20622 12832 20628 12844
rect 19935 12804 20628 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 13722 12764 13728 12776
rect 13412 12736 13584 12764
rect 13683 12736 13728 12764
rect 13412 12724 13418 12736
rect 13722 12724 13728 12736
rect 13780 12764 13786 12776
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 13780 12736 16129 12764
rect 13780 12724 13786 12736
rect 16117 12733 16129 12736
rect 16163 12764 16175 12767
rect 16206 12764 16212 12776
rect 16163 12736 16212 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 18138 12764 18144 12776
rect 16724 12736 18144 12764
rect 16724 12724 16730 12736
rect 18138 12724 18144 12736
rect 18196 12764 18202 12776
rect 18432 12764 18460 12795
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 22002 12832 22008 12844
rect 20763 12804 22008 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22554 12832 22560 12844
rect 22327 12804 22560 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22554 12792 22560 12804
rect 22612 12792 22618 12844
rect 18196 12736 18460 12764
rect 18196 12724 18202 12736
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20312 12736 20453 12764
rect 20312 12724 20318 12736
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 20441 12727 20499 12733
rect 20901 12767 20959 12773
rect 20901 12733 20913 12767
rect 20947 12733 20959 12767
rect 22370 12764 22376 12776
rect 22331 12736 22376 12764
rect 20901 12727 20959 12733
rect 14274 12696 14280 12708
rect 13188 12668 14280 12696
rect 14274 12656 14280 12668
rect 14332 12696 14338 12708
rect 16853 12699 16911 12705
rect 16853 12696 16865 12699
rect 14332 12668 16865 12696
rect 14332 12656 14338 12668
rect 16853 12665 16865 12668
rect 16899 12665 16911 12699
rect 16853 12659 16911 12665
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 13354 12628 13360 12640
rect 12115 12600 13360 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 14366 12628 14372 12640
rect 13504 12600 14372 12628
rect 13504 12588 13510 12600
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 14826 12628 14832 12640
rect 14739 12600 14832 12628
rect 14826 12588 14832 12600
rect 14884 12628 14890 12640
rect 15838 12628 15844 12640
rect 14884 12600 15844 12628
rect 14884 12588 14890 12600
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17184 12600 17509 12628
rect 17184 12588 17190 12600
rect 17497 12597 17509 12600
rect 17543 12628 17555 12631
rect 20162 12628 20168 12640
rect 17543 12600 20168 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 20162 12588 20168 12600
rect 20220 12628 20226 12640
rect 20916 12628 20944 12727
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 23750 12656 23756 12708
rect 23808 12696 23814 12708
rect 25317 12699 25375 12705
rect 25317 12696 25329 12699
rect 23808 12668 25329 12696
rect 23808 12656 23814 12668
rect 25317 12665 25329 12668
rect 25363 12665 25375 12699
rect 25317 12659 25375 12665
rect 21082 12628 21088 12640
rect 20220 12600 21088 12628
rect 20220 12588 20226 12600
rect 21082 12588 21088 12600
rect 21140 12628 21146 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 21140 12600 21189 12628
rect 21140 12588 21146 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 23198 12628 23204 12640
rect 23159 12600 23204 12628
rect 21177 12591 21235 12597
rect 23198 12588 23204 12600
rect 23256 12588 23262 12640
rect 1104 12538 28336 12560
rect 1104 12486 3282 12538
rect 3334 12486 3346 12538
rect 3398 12486 3410 12538
rect 3462 12486 3474 12538
rect 3526 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 6410 12538
rect 6462 12486 6474 12538
rect 6526 12486 9282 12538
rect 9334 12486 9346 12538
rect 9398 12486 9410 12538
rect 9462 12486 9474 12538
rect 9526 12486 12282 12538
rect 12334 12486 12346 12538
rect 12398 12486 12410 12538
rect 12462 12486 12474 12538
rect 12526 12486 15282 12538
rect 15334 12486 15346 12538
rect 15398 12486 15410 12538
rect 15462 12486 15474 12538
rect 15526 12486 18282 12538
rect 18334 12486 18346 12538
rect 18398 12486 18410 12538
rect 18462 12486 18474 12538
rect 18526 12486 21282 12538
rect 21334 12486 21346 12538
rect 21398 12486 21410 12538
rect 21462 12486 21474 12538
rect 21526 12486 24282 12538
rect 24334 12486 24346 12538
rect 24398 12486 24410 12538
rect 24462 12486 24474 12538
rect 24526 12486 27282 12538
rect 27334 12486 27346 12538
rect 27398 12486 27410 12538
rect 27462 12486 27474 12538
rect 27526 12486 28336 12538
rect 1104 12464 28336 12486
rect 9122 12424 9128 12436
rect 9083 12396 9128 12424
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12424 11299 12427
rect 11514 12424 11520 12436
rect 11287 12396 11520 12424
rect 11287 12393 11299 12396
rect 11241 12387 11299 12393
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 13817 12427 13875 12433
rect 13817 12424 13829 12427
rect 13688 12396 13829 12424
rect 13688 12384 13694 12396
rect 13817 12393 13829 12396
rect 13863 12393 13875 12427
rect 14274 12424 14280 12436
rect 14235 12396 14280 12424
rect 13817 12387 13875 12393
rect 14274 12384 14280 12396
rect 14332 12384 14338 12436
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 16724 12396 17049 12424
rect 16724 12384 16730 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 17678 12424 17684 12436
rect 17639 12396 17684 12424
rect 17037 12387 17095 12393
rect 15930 12356 15936 12368
rect 15891 12328 15936 12356
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 8202 12288 8208 12300
rect 8115 12260 8208 12288
rect 8202 12248 8208 12260
rect 8260 12288 8266 12300
rect 8662 12288 8668 12300
rect 8260 12260 8668 12288
rect 8260 12248 8266 12260
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 11790 12288 11796 12300
rect 11751 12260 11796 12288
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12288 15531 12291
rect 15838 12288 15844 12300
rect 15519 12260 15844 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 17052 12288 17080 12387
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 19061 12427 19119 12433
rect 19061 12424 19073 12427
rect 17828 12396 19073 12424
rect 17828 12384 17834 12396
rect 19061 12393 19073 12396
rect 19107 12393 19119 12427
rect 20254 12424 20260 12436
rect 20215 12396 20260 12424
rect 19061 12387 19119 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 23198 12384 23204 12436
rect 23256 12424 23262 12436
rect 24397 12427 24455 12433
rect 24397 12424 24409 12427
rect 23256 12396 24409 12424
rect 23256 12384 23262 12396
rect 24397 12393 24409 12396
rect 24443 12393 24455 12427
rect 24397 12387 24455 12393
rect 18325 12359 18383 12365
rect 18325 12325 18337 12359
rect 18371 12356 18383 12359
rect 18598 12356 18604 12368
rect 18371 12328 18604 12356
rect 18371 12325 18383 12328
rect 18325 12319 18383 12325
rect 17405 12291 17463 12297
rect 17405 12288 17417 12291
rect 17052 12260 17417 12288
rect 17405 12257 17417 12260
rect 17451 12257 17463 12291
rect 17405 12251 17463 12257
rect 8294 12220 8300 12232
rect 8255 12192 8300 12220
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11480 12192 11529 12220
rect 11480 12180 11486 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 16206 12220 16212 12232
rect 16167 12192 16212 12220
rect 11517 12183 11575 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 16482 12220 16488 12232
rect 16443 12192 16488 12220
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 17310 12180 17316 12232
rect 17368 12220 17374 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 17368 12192 17509 12220
rect 17368 12180 17374 12192
rect 17497 12189 17509 12192
rect 17543 12220 17555 12223
rect 18340 12220 18368 12319
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 18748 12328 21281 12356
rect 18748 12316 18754 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 22189 12359 22247 12365
rect 22189 12325 22201 12359
rect 22235 12356 22247 12359
rect 22646 12356 22652 12368
rect 22235 12328 22652 12356
rect 22235 12325 22247 12328
rect 22189 12319 22247 12325
rect 22646 12316 22652 12328
rect 22704 12316 22710 12368
rect 25133 12359 25191 12365
rect 25133 12325 25145 12359
rect 25179 12356 25191 12359
rect 28718 12356 28724 12368
rect 25179 12328 28724 12356
rect 25179 12325 25191 12328
rect 25133 12319 25191 12325
rect 28718 12316 28724 12328
rect 28776 12316 28782 12368
rect 17543 12192 18368 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 18969 12223 19027 12229
rect 18969 12220 18981 12223
rect 18932 12192 18981 12220
rect 18932 12180 18938 12192
rect 18969 12189 18981 12192
rect 19015 12189 19027 12223
rect 21082 12220 21088 12232
rect 21043 12192 21088 12220
rect 18969 12183 19027 12189
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 22370 12220 22376 12232
rect 22331 12192 22376 12220
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22554 12220 22560 12232
rect 22515 12192 22560 12220
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 22741 12223 22799 12229
rect 22741 12220 22753 12223
rect 22704 12192 22753 12220
rect 22704 12180 22710 12192
rect 22741 12189 22753 12192
rect 22787 12220 22799 12223
rect 23750 12220 23756 12232
rect 22787 12192 23756 12220
rect 22787 12189 22799 12192
rect 22741 12183 22799 12189
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 8757 12155 8815 12161
rect 8757 12121 8769 12155
rect 8803 12152 8815 12155
rect 9858 12152 9864 12164
rect 8803 12124 9864 12152
rect 8803 12121 8815 12124
rect 8757 12115 8815 12121
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 12250 12112 12256 12164
rect 12308 12112 12314 12164
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12152 13599 12155
rect 13722 12152 13728 12164
rect 13587 12124 13728 12152
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 10873 12087 10931 12093
rect 10873 12053 10885 12087
rect 10919 12084 10931 12087
rect 12802 12084 12808 12096
rect 10919 12056 12808 12084
rect 10919 12053 10931 12056
rect 10873 12047 10931 12053
rect 12802 12044 12808 12056
rect 12860 12084 12866 12096
rect 13556 12084 13584 12115
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 18782 12152 18788 12164
rect 18743 12124 18788 12152
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 22572 12152 22600 12180
rect 23201 12155 23259 12161
rect 23201 12152 23213 12155
rect 22572 12124 23213 12152
rect 23201 12121 23213 12124
rect 23247 12121 23259 12155
rect 23201 12115 23259 12121
rect 12860 12056 13584 12084
rect 14921 12087 14979 12093
rect 12860 12044 12866 12056
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15102 12084 15108 12096
rect 14967 12056 15108 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 19981 12087 20039 12093
rect 19981 12053 19993 12087
rect 20027 12084 20039 12087
rect 20162 12084 20168 12096
rect 20027 12056 20168 12084
rect 20027 12053 20039 12056
rect 19981 12047 20039 12053
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 21637 12087 21695 12093
rect 21637 12053 21649 12087
rect 21683 12084 21695 12087
rect 22002 12084 22008 12096
rect 21683 12056 22008 12084
rect 21683 12053 21695 12056
rect 21637 12047 21695 12053
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 1104 11994 28336 12016
rect 1104 11942 1782 11994
rect 1834 11942 1846 11994
rect 1898 11942 1910 11994
rect 1962 11942 1974 11994
rect 2026 11942 4782 11994
rect 4834 11942 4846 11994
rect 4898 11942 4910 11994
rect 4962 11942 4974 11994
rect 5026 11942 7782 11994
rect 7834 11942 7846 11994
rect 7898 11942 7910 11994
rect 7962 11942 7974 11994
rect 8026 11942 10782 11994
rect 10834 11942 10846 11994
rect 10898 11942 10910 11994
rect 10962 11942 10974 11994
rect 11026 11942 13782 11994
rect 13834 11942 13846 11994
rect 13898 11942 13910 11994
rect 13962 11942 13974 11994
rect 14026 11942 16782 11994
rect 16834 11942 16846 11994
rect 16898 11942 16910 11994
rect 16962 11942 16974 11994
rect 17026 11942 19782 11994
rect 19834 11942 19846 11994
rect 19898 11942 19910 11994
rect 19962 11942 19974 11994
rect 20026 11942 22782 11994
rect 22834 11942 22846 11994
rect 22898 11942 22910 11994
rect 22962 11942 22974 11994
rect 23026 11942 25782 11994
rect 25834 11942 25846 11994
rect 25898 11942 25910 11994
rect 25962 11942 25974 11994
rect 26026 11942 28336 11994
rect 1104 11920 28336 11942
rect 8202 11880 8208 11892
rect 8163 11852 8208 11880
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8352 11852 8585 11880
rect 8352 11840 8358 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 10735 11852 11529 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 11517 11849 11529 11852
rect 11563 11880 11575 11883
rect 12250 11880 12256 11892
rect 11563 11852 12256 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 13262 11880 13268 11892
rect 13219 11852 13268 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13596 11852 13645 11880
rect 13596 11840 13602 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14550 11880 14556 11892
rect 14139 11852 14556 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 16574 11880 16580 11892
rect 16535 11852 16580 11880
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17368 11852 17417 11880
rect 17368 11840 17374 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 18138 11840 18144 11892
rect 18196 11880 18202 11892
rect 18233 11883 18291 11889
rect 18233 11880 18245 11883
rect 18196 11852 18245 11880
rect 18196 11840 18202 11852
rect 18233 11849 18245 11852
rect 18279 11849 18291 11883
rect 18233 11843 18291 11849
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 20441 11883 20499 11889
rect 20441 11880 20453 11883
rect 18840 11852 20453 11880
rect 18840 11840 18846 11852
rect 20441 11849 20453 11852
rect 20487 11849 20499 11883
rect 20441 11843 20499 11849
rect 22370 11840 22376 11892
rect 22428 11880 22434 11892
rect 22741 11883 22799 11889
rect 22741 11880 22753 11883
rect 22428 11852 22753 11880
rect 22428 11840 22434 11852
rect 22741 11849 22753 11852
rect 22787 11849 22799 11883
rect 22741 11843 22799 11849
rect 11057 11815 11115 11821
rect 11057 11781 11069 11815
rect 11103 11812 11115 11815
rect 11790 11812 11796 11824
rect 11103 11784 11796 11812
rect 11103 11781 11115 11784
rect 11057 11775 11115 11781
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 14274 11772 14280 11824
rect 14332 11812 14338 11824
rect 20714 11812 20720 11824
rect 14332 11784 15240 11812
rect 14332 11772 14338 11784
rect 9766 11744 9772 11756
rect 9727 11716 9772 11744
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 11333 11747 11391 11753
rect 9876 11716 11284 11744
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11676 8999 11679
rect 9122 11676 9128 11688
rect 8987 11648 9128 11676
rect 8987 11645 8999 11648
rect 8941 11639 8999 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9582 11676 9588 11688
rect 9539 11648 9588 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9582 11636 9588 11648
rect 9640 11676 9646 11688
rect 9876 11676 9904 11716
rect 9640 11648 9904 11676
rect 9953 11679 10011 11685
rect 9640 11636 9646 11648
rect 9953 11645 9965 11679
rect 9999 11645 10011 11679
rect 11256 11676 11284 11716
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11514 11744 11520 11756
rect 11379 11716 11520 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 12618 11744 12624 11756
rect 11624 11716 12624 11744
rect 11624 11676 11652 11716
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 14918 11744 14924 11756
rect 14879 11716 14924 11744
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15212 11753 15240 11784
rect 18984 11784 20720 11812
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16482 11744 16488 11756
rect 15887 11716 16488 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11744 17003 11747
rect 17126 11744 17132 11756
rect 16991 11716 17132 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 18984 11753 19012 11784
rect 20714 11772 20720 11784
rect 20772 11772 20778 11824
rect 20990 11812 20996 11824
rect 20951 11784 20996 11812
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 21082 11772 21088 11824
rect 21140 11812 21146 11824
rect 23109 11815 23167 11821
rect 23109 11812 23121 11815
rect 21140 11784 23121 11812
rect 21140 11772 21146 11784
rect 23109 11781 23121 11784
rect 23155 11781 23167 11815
rect 23109 11775 23167 11781
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 19426 11744 19432 11756
rect 19387 11716 19432 11744
rect 18969 11707 19027 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 19702 11744 19708 11756
rect 19567 11716 19708 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 19702 11704 19708 11716
rect 19760 11744 19766 11756
rect 20254 11744 20260 11756
rect 19760 11716 20260 11744
rect 19760 11704 19766 11716
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 21100 11744 21128 11772
rect 20496 11716 21128 11744
rect 21729 11747 21787 11753
rect 20496 11704 20502 11716
rect 21729 11713 21741 11747
rect 21775 11744 21787 11747
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 21775 11716 22385 11744
rect 21775 11713 21787 11716
rect 21729 11707 21787 11713
rect 22373 11713 22385 11716
rect 22419 11744 22431 11747
rect 22554 11744 22560 11756
rect 22419 11716 22560 11744
rect 22419 11713 22431 11716
rect 22373 11707 22431 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 11256 11648 11652 11676
rect 9953 11639 10011 11645
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 9968 11608 9996 11639
rect 14090 11636 14096 11688
rect 14148 11676 14154 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14148 11648 14381 11676
rect 14148 11636 14154 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 15654 11676 15660 11688
rect 15615 11648 15660 11676
rect 14369 11639 14427 11645
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 18598 11636 18604 11688
rect 18656 11676 18662 11688
rect 18785 11679 18843 11685
rect 18785 11676 18797 11679
rect 18656 11648 18797 11676
rect 18656 11636 18662 11648
rect 18785 11645 18797 11648
rect 18831 11645 18843 11679
rect 18785 11639 18843 11645
rect 21082 11636 21088 11688
rect 21140 11676 21146 11688
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21140 11648 21373 11676
rect 21140 11636 21146 11648
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 8628 11580 9996 11608
rect 8628 11568 8634 11580
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 11664 11580 12817 11608
rect 11664 11568 11670 11580
rect 12805 11577 12817 11580
rect 12851 11608 12863 11611
rect 13170 11608 13176 11620
rect 12851 11580 13176 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 21269 11611 21327 11617
rect 21269 11608 21281 11611
rect 19996 11580 21281 11608
rect 19996 11552 20024 11580
rect 21269 11577 21281 11580
rect 21315 11577 21327 11611
rect 21269 11571 21327 11577
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11480 11512 11805 11540
rect 11480 11500 11486 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 16209 11543 16267 11549
rect 16209 11509 16221 11543
rect 16255 11540 16267 11543
rect 16298 11540 16304 11552
rect 16255 11512 16304 11540
rect 16255 11509 16267 11512
rect 16209 11503 16267 11509
rect 16298 11500 16304 11512
rect 16356 11540 16362 11552
rect 16666 11540 16672 11552
rect 16356 11512 16672 11540
rect 16356 11500 16362 11512
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 19978 11540 19984 11552
rect 19939 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 21131 11543 21189 11549
rect 21131 11540 21143 11543
rect 20680 11512 21143 11540
rect 20680 11500 20686 11512
rect 21131 11509 21143 11512
rect 21177 11540 21189 11543
rect 21818 11540 21824 11552
rect 21177 11512 21824 11540
rect 21177 11509 21189 11512
rect 21131 11503 21189 11509
rect 21818 11500 21824 11512
rect 21876 11500 21882 11552
rect 22002 11540 22008 11552
rect 21963 11512 22008 11540
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 1104 11450 28336 11472
rect 1104 11398 3282 11450
rect 3334 11398 3346 11450
rect 3398 11398 3410 11450
rect 3462 11398 3474 11450
rect 3526 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 6410 11450
rect 6462 11398 6474 11450
rect 6526 11398 9282 11450
rect 9334 11398 9346 11450
rect 9398 11398 9410 11450
rect 9462 11398 9474 11450
rect 9526 11398 12282 11450
rect 12334 11398 12346 11450
rect 12398 11398 12410 11450
rect 12462 11398 12474 11450
rect 12526 11398 15282 11450
rect 15334 11398 15346 11450
rect 15398 11398 15410 11450
rect 15462 11398 15474 11450
rect 15526 11398 18282 11450
rect 18334 11398 18346 11450
rect 18398 11398 18410 11450
rect 18462 11398 18474 11450
rect 18526 11398 21282 11450
rect 21334 11398 21346 11450
rect 21398 11398 21410 11450
rect 21462 11398 21474 11450
rect 21526 11398 24282 11450
rect 24334 11398 24346 11450
rect 24398 11398 24410 11450
rect 24462 11398 24474 11450
rect 24526 11398 27282 11450
rect 27334 11398 27346 11450
rect 27398 11398 27410 11450
rect 27462 11398 27474 11450
rect 27526 11398 28336 11450
rect 1104 11376 28336 11398
rect 8665 11339 8723 11345
rect 8665 11305 8677 11339
rect 8711 11336 8723 11339
rect 9766 11336 9772 11348
rect 8711 11308 9772 11336
rect 8711 11305 8723 11308
rect 8665 11299 8723 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12860 11308 12909 11336
rect 12860 11296 12866 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 12897 11299 12955 11305
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13228 11308 13277 11336
rect 13228 11296 13234 11308
rect 13265 11305 13277 11308
rect 13311 11336 13323 11339
rect 13725 11339 13783 11345
rect 13311 11308 13584 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 9582 11268 9588 11280
rect 9079 11240 9588 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 11388 11172 12081 11200
rect 11388 11160 11394 11172
rect 12069 11169 12081 11172
rect 12115 11200 12127 11203
rect 13262 11200 13268 11212
rect 12115 11172 13268 11200
rect 12115 11169 12127 11172
rect 12069 11163 12127 11169
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 11241 11135 11299 11141
rect 11241 11101 11253 11135
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 11606 11132 11612 11144
rect 11567 11104 11612 11132
rect 11425 11095 11483 11101
rect 10781 11067 10839 11073
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 11146 11064 11152 11076
rect 10827 11036 11152 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 8297 10999 8355 11005
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 8570 10996 8576 11008
rect 8343 10968 8576 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 10410 10996 10416 11008
rect 10371 10968 10416 10996
rect 10410 10956 10416 10968
rect 10468 10996 10474 11008
rect 11256 10996 11284 11095
rect 10468 10968 11284 10996
rect 11440 10996 11468 11095
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 12158 11132 12164 11144
rect 12119 11104 12164 11132
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 13556 11132 13584 11308
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 14918 11336 14924 11348
rect 13771 11308 14924 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 14918 11296 14924 11308
rect 14976 11336 14982 11348
rect 15565 11339 15623 11345
rect 15565 11336 15577 11339
rect 14976 11308 15577 11336
rect 14976 11296 14982 11308
rect 15565 11305 15577 11308
rect 15611 11305 15623 11339
rect 15565 11299 15623 11305
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 19702 11336 19708 11348
rect 16540 11308 18276 11336
rect 19663 11308 19708 11336
rect 16540 11296 16546 11308
rect 13630 11228 13636 11280
rect 13688 11268 13694 11280
rect 14274 11268 14280 11280
rect 13688 11240 14280 11268
rect 13688 11228 13694 11240
rect 14274 11228 14280 11240
rect 14332 11228 14338 11280
rect 14826 11268 14832 11280
rect 14787 11240 14832 11268
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 16264 11240 16712 11268
rect 16264 11228 16270 11240
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 16022 11200 16028 11212
rect 14424 11172 16028 11200
rect 14424 11160 14430 11172
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 16448 11172 16589 11200
rect 16448 11160 16454 11172
rect 16577 11169 16589 11172
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 15654 11132 15660 11144
rect 13556 11104 15660 11132
rect 15654 11092 15660 11104
rect 15712 11092 15718 11144
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 15988 11104 16129 11132
rect 15988 11092 15994 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 16117 11095 16175 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16684 11132 16712 11240
rect 18248 11209 18276 11308
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 20036 11308 20453 11336
rect 20036 11296 20042 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 22002 11336 22008 11348
rect 21963 11308 22008 11336
rect 20441 11299 20499 11305
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22646 11296 22652 11348
rect 22704 11336 22710 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22704 11308 22937 11336
rect 22704 11296 22710 11308
rect 22925 11305 22937 11308
rect 22971 11305 22983 11339
rect 22925 11299 22983 11305
rect 21818 11228 21824 11280
rect 21876 11268 21882 11280
rect 22557 11271 22615 11277
rect 22557 11268 22569 11271
rect 21876 11240 22569 11268
rect 21876 11228 21882 11240
rect 22557 11237 22569 11240
rect 22603 11237 22615 11271
rect 22557 11231 22615 11237
rect 18233 11203 18291 11209
rect 18233 11169 18245 11203
rect 18279 11200 18291 11203
rect 22462 11200 22468 11212
rect 18279 11172 22468 11200
rect 18279 11169 18291 11172
rect 18233 11163 18291 11169
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 16684 11104 17785 11132
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 14093 11067 14151 11073
rect 14093 11033 14105 11067
rect 14139 11064 14151 11067
rect 15102 11064 15108 11076
rect 14139 11036 15108 11064
rect 14139 11033 14151 11036
rect 14093 11027 14151 11033
rect 15102 11024 15108 11036
rect 15160 11064 15166 11076
rect 17313 11067 17371 11073
rect 17313 11064 17325 11067
rect 15160 11036 17325 11064
rect 15160 11024 15166 11036
rect 17313 11033 17325 11036
rect 17359 11033 17371 11067
rect 17313 11027 17371 11033
rect 18156 11064 18184 11095
rect 19242 11092 19248 11144
rect 19300 11132 19306 11144
rect 19337 11135 19395 11141
rect 19337 11132 19349 11135
rect 19300 11104 19349 11132
rect 19300 11092 19306 11104
rect 19337 11101 19349 11104
rect 19383 11101 19395 11135
rect 21634 11132 21640 11144
rect 21595 11104 21640 11132
rect 19337 11095 19395 11101
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 19426 11064 19432 11076
rect 18156 11036 19432 11064
rect 11882 10996 11888 11008
rect 11440 10968 11888 10996
rect 10468 10956 10474 10968
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 11974 10956 11980 11008
rect 12032 10996 12038 11008
rect 12529 10999 12587 11005
rect 12529 10996 12541 10999
rect 12032 10968 12541 10996
rect 12032 10956 12038 10968
rect 12529 10965 12541 10968
rect 12575 10996 12587 10999
rect 12618 10996 12624 11008
rect 12575 10968 12624 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 14332 10968 14381 10996
rect 14332 10956 14338 10968
rect 14369 10965 14381 10968
rect 14415 10965 14427 10999
rect 14369 10959 14427 10965
rect 17037 10999 17095 11005
rect 17037 10965 17049 10999
rect 17083 10996 17095 10999
rect 17126 10996 17132 11008
rect 17083 10968 17132 10996
rect 17083 10965 17095 10968
rect 17037 10959 17095 10965
rect 17126 10956 17132 10968
rect 17184 10996 17190 11008
rect 18156 10996 18184 11036
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 17184 10968 18184 10996
rect 17184 10956 17190 10968
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 18785 10999 18843 11005
rect 18785 10996 18797 10999
rect 18656 10968 18797 10996
rect 18656 10956 18662 10968
rect 18785 10965 18797 10968
rect 18831 10965 18843 10999
rect 21082 10996 21088 11008
rect 21043 10968 21088 10996
rect 18785 10959 18843 10965
rect 21082 10956 21088 10968
rect 21140 10956 21146 11008
rect 1104 10906 28336 10928
rect 1104 10854 1782 10906
rect 1834 10854 1846 10906
rect 1898 10854 1910 10906
rect 1962 10854 1974 10906
rect 2026 10854 4782 10906
rect 4834 10854 4846 10906
rect 4898 10854 4910 10906
rect 4962 10854 4974 10906
rect 5026 10854 7782 10906
rect 7834 10854 7846 10906
rect 7898 10854 7910 10906
rect 7962 10854 7974 10906
rect 8026 10854 10782 10906
rect 10834 10854 10846 10906
rect 10898 10854 10910 10906
rect 10962 10854 10974 10906
rect 11026 10854 13782 10906
rect 13834 10854 13846 10906
rect 13898 10854 13910 10906
rect 13962 10854 13974 10906
rect 14026 10854 16782 10906
rect 16834 10854 16846 10906
rect 16898 10854 16910 10906
rect 16962 10854 16974 10906
rect 17026 10854 19782 10906
rect 19834 10854 19846 10906
rect 19898 10854 19910 10906
rect 19962 10854 19974 10906
rect 20026 10854 22782 10906
rect 22834 10854 22846 10906
rect 22898 10854 22910 10906
rect 22962 10854 22974 10906
rect 23026 10854 25782 10906
rect 25834 10854 25846 10906
rect 25898 10854 25910 10906
rect 25962 10854 25974 10906
rect 26026 10854 28336 10906
rect 1104 10832 28336 10854
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9769 10795 9827 10801
rect 8352 10764 9352 10792
rect 8352 10752 8358 10764
rect 8662 10684 8668 10736
rect 8720 10724 8726 10736
rect 9030 10724 9036 10736
rect 8720 10696 9036 10724
rect 8720 10684 8726 10696
rect 9030 10684 9036 10696
rect 9088 10724 9094 10736
rect 9088 10696 9260 10724
rect 9088 10684 9094 10696
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10656 7711 10659
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 7699 10628 8309 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 8297 10625 8309 10628
rect 8343 10656 8355 10659
rect 8754 10656 8760 10668
rect 8343 10628 8760 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9232 10665 9260 10696
rect 9324 10665 9352 10764
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 9815 10764 11253 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 11241 10761 11253 10764
rect 11287 10792 11299 10795
rect 12158 10792 12164 10804
rect 11287 10764 12164 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 13081 10795 13139 10801
rect 13081 10792 13093 10795
rect 12759 10764 13093 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 13081 10761 13093 10764
rect 13127 10792 13139 10795
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 13127 10764 13461 10792
rect 13127 10761 13139 10764
rect 13081 10755 13139 10761
rect 13449 10761 13461 10764
rect 13495 10792 13507 10795
rect 16022 10792 16028 10804
rect 13495 10764 15792 10792
rect 15983 10764 16028 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 10873 10727 10931 10733
rect 10873 10693 10885 10727
rect 10919 10724 10931 10727
rect 11330 10724 11336 10736
rect 10919 10696 11336 10724
rect 10919 10693 10931 10696
rect 10873 10687 10931 10693
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 10318 10656 10324 10668
rect 9355 10628 10324 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8202 10588 8208 10600
rect 7791 10560 8208 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 10888 10520 10916 10687
rect 11330 10684 11336 10696
rect 11388 10724 11394 10736
rect 11698 10724 11704 10736
rect 11388 10696 11704 10724
rect 11388 10684 11394 10696
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 14458 10684 14464 10736
rect 14516 10684 14522 10736
rect 15764 10733 15792 10764
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 19337 10795 19395 10801
rect 19337 10792 19349 10795
rect 17543 10764 19349 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10724 15807 10727
rect 16482 10724 16488 10736
rect 15795 10696 16488 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 18984 10733 19012 10764
rect 19337 10761 19349 10764
rect 19383 10792 19395 10795
rect 19426 10792 19432 10804
rect 19383 10764 19432 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19610 10792 19616 10804
rect 19571 10764 19616 10792
rect 19610 10752 19616 10764
rect 19668 10752 19674 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 20772 10764 22017 10792
rect 20772 10752 20778 10764
rect 18969 10727 19027 10733
rect 18969 10693 18981 10727
rect 19015 10693 19027 10727
rect 18969 10687 19027 10693
rect 20165 10727 20223 10733
rect 20165 10693 20177 10727
rect 20211 10724 20223 10727
rect 21082 10724 21088 10736
rect 20211 10696 21088 10724
rect 20211 10693 20223 10696
rect 20165 10687 20223 10693
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 11514 10656 11520 10668
rect 11475 10628 11520 10656
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 15654 10616 15660 10668
rect 15712 10656 15718 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 15712 10628 16957 10656
rect 15712 10616 15718 10628
rect 16945 10625 16957 10628
rect 16991 10656 17003 10659
rect 17586 10656 17592 10668
rect 16991 10628 17592 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 17586 10616 17592 10628
rect 17644 10616 17650 10668
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 19150 10656 19156 10668
rect 18923 10628 19156 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 19150 10616 19156 10628
rect 19208 10656 19214 10668
rect 20438 10656 20444 10668
rect 19208 10628 20444 10656
rect 19208 10616 19214 10628
rect 20438 10616 20444 10628
rect 20496 10616 20502 10668
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 21284 10665 21312 10764
rect 22005 10761 22017 10764
rect 22051 10792 22063 10795
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22051 10764 22385 10792
rect 22051 10761 22063 10764
rect 22005 10755 22063 10761
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22741 10795 22799 10801
rect 22741 10792 22753 10795
rect 22520 10764 22753 10792
rect 22520 10752 22526 10764
rect 22741 10761 22753 10764
rect 22787 10761 22799 10795
rect 22741 10755 22799 10761
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 13538 10548 13544 10600
rect 13596 10588 13602 10600
rect 13725 10591 13783 10597
rect 13725 10588 13737 10591
rect 13596 10560 13737 10588
rect 13596 10548 13602 10560
rect 13725 10557 13737 10560
rect 13771 10557 13783 10591
rect 13998 10588 14004 10600
rect 13959 10560 14004 10588
rect 13725 10551 13783 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 20346 10548 20352 10600
rect 20404 10588 20410 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20404 10560 20729 10588
rect 20404 10548 20410 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 21192 10532 21220 10619
rect 9646 10492 10916 10520
rect 16669 10523 16727 10529
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 8846 10452 8852 10464
rect 8628 10424 8852 10452
rect 8628 10412 8634 10424
rect 8846 10412 8852 10424
rect 8904 10452 8910 10464
rect 9646 10452 9674 10492
rect 16669 10489 16681 10523
rect 16715 10520 16727 10523
rect 19242 10520 19248 10532
rect 16715 10492 19248 10520
rect 16715 10489 16727 10492
rect 16669 10483 16727 10489
rect 19242 10480 19248 10492
rect 19300 10520 19306 10532
rect 21174 10520 21180 10532
rect 19300 10492 21180 10520
rect 19300 10480 19306 10492
rect 21174 10480 21180 10492
rect 21232 10480 21238 10532
rect 22002 10520 22008 10532
rect 21376 10492 22008 10520
rect 8904 10424 9674 10452
rect 10505 10455 10563 10461
rect 8904 10412 8910 10424
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 11606 10452 11612 10464
rect 10551 10424 11612 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 11882 10452 11888 10464
rect 11843 10424 11888 10452
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 16758 10412 16764 10464
rect 16816 10452 16822 10464
rect 17129 10455 17187 10461
rect 17129 10452 17141 10455
rect 16816 10424 17141 10452
rect 16816 10412 16822 10424
rect 17129 10421 17141 10424
rect 17175 10452 17187 10455
rect 17954 10452 17960 10464
rect 17175 10424 17960 10452
rect 17175 10421 17187 10424
rect 17129 10415 17187 10421
rect 17954 10412 17960 10424
rect 18012 10452 18018 10464
rect 21376 10452 21404 10492
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 21634 10452 21640 10464
rect 18012 10424 21404 10452
rect 21595 10424 21640 10452
rect 18012 10412 18018 10424
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 1104 10362 28336 10384
rect 1104 10310 3282 10362
rect 3334 10310 3346 10362
rect 3398 10310 3410 10362
rect 3462 10310 3474 10362
rect 3526 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 6410 10362
rect 6462 10310 6474 10362
rect 6526 10310 9282 10362
rect 9334 10310 9346 10362
rect 9398 10310 9410 10362
rect 9462 10310 9474 10362
rect 9526 10310 12282 10362
rect 12334 10310 12346 10362
rect 12398 10310 12410 10362
rect 12462 10310 12474 10362
rect 12526 10310 15282 10362
rect 15334 10310 15346 10362
rect 15398 10310 15410 10362
rect 15462 10310 15474 10362
rect 15526 10310 18282 10362
rect 18334 10310 18346 10362
rect 18398 10310 18410 10362
rect 18462 10310 18474 10362
rect 18526 10310 21282 10362
rect 21334 10310 21346 10362
rect 21398 10310 21410 10362
rect 21462 10310 21474 10362
rect 21526 10310 24282 10362
rect 24334 10310 24346 10362
rect 24398 10310 24410 10362
rect 24462 10310 24474 10362
rect 24526 10310 27282 10362
rect 27334 10310 27346 10362
rect 27398 10310 27410 10362
rect 27462 10310 27474 10362
rect 27526 10310 28336 10362
rect 1104 10288 28336 10310
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 8754 10248 8760 10260
rect 6503 10220 8760 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 8754 10208 8760 10220
rect 8812 10248 8818 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 8812 10220 10057 10248
rect 8812 10208 8818 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 10045 10211 10103 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 14056 10220 14565 10248
rect 14056 10208 14062 10220
rect 14553 10217 14565 10220
rect 14599 10217 14611 10251
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 14553 10211 14611 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 20070 10248 20076 10260
rect 19015 10220 20076 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20346 10248 20352 10260
rect 20307 10220 20352 10248
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20990 10208 20996 10260
rect 21048 10248 21054 10260
rect 21085 10251 21143 10257
rect 21085 10248 21097 10251
rect 21048 10220 21097 10248
rect 21048 10208 21054 10220
rect 21085 10217 21097 10220
rect 21131 10217 21143 10251
rect 21085 10211 21143 10217
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21453 10251 21511 10257
rect 21453 10248 21465 10251
rect 21232 10220 21465 10248
rect 21232 10208 21238 10220
rect 21453 10217 21465 10220
rect 21499 10217 21511 10251
rect 21453 10211 21511 10217
rect 9030 10180 9036 10192
rect 8991 10152 9036 10180
rect 9030 10140 9036 10152
rect 9088 10140 9094 10192
rect 13449 10183 13507 10189
rect 13449 10149 13461 10183
rect 13495 10180 13507 10183
rect 13909 10183 13967 10189
rect 13909 10180 13921 10183
rect 13495 10152 13921 10180
rect 13495 10149 13507 10152
rect 13449 10143 13507 10149
rect 13909 10149 13921 10152
rect 13955 10180 13967 10183
rect 14458 10180 14464 10192
rect 13955 10152 14464 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 15565 10183 15623 10189
rect 15565 10149 15577 10183
rect 15611 10180 15623 10183
rect 16390 10180 16396 10192
rect 15611 10152 16396 10180
rect 15611 10149 15623 10152
rect 15565 10143 15623 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 19521 10183 19579 10189
rect 19521 10180 19533 10183
rect 18984 10152 19533 10180
rect 18984 10124 19012 10152
rect 19521 10149 19533 10152
rect 19567 10149 19579 10183
rect 19521 10143 19579 10149
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7098 10112 7104 10124
rect 6779 10084 7104 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 11146 10112 11152 10124
rect 11107 10084 11152 10112
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 11572 10084 13124 10112
rect 11572 10072 11578 10084
rect 9858 10044 9864 10056
rect 9819 10016 9864 10044
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10013 10931 10047
rect 13096 10044 13124 10084
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15712 10084 16712 10112
rect 15712 10072 15718 10084
rect 13630 10044 13636 10056
rect 13096 10016 13636 10044
rect 10873 10007 10931 10013
rect 7006 9976 7012 9988
rect 6967 9948 7012 9976
rect 7006 9936 7012 9948
rect 7064 9936 7070 9988
rect 7466 9936 7472 9988
rect 7524 9936 7530 9988
rect 8754 9976 8760 9988
rect 8715 9948 8760 9976
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 10888 9976 10916 10007
rect 13630 10004 13636 10016
rect 13688 10044 13694 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13688 10016 13737 10044
rect 13688 10004 13694 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 16574 10044 16580 10056
rect 16535 10016 16580 10044
rect 13725 10007 13783 10013
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 16684 10053 16712 10084
rect 18966 10072 18972 10124
rect 19024 10072 19030 10124
rect 19610 10112 19616 10124
rect 19523 10084 19616 10112
rect 19610 10072 19616 10084
rect 19668 10112 19674 10124
rect 20364 10112 20392 10208
rect 19668 10084 20392 10112
rect 19668 10072 19674 10084
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10044 16727 10047
rect 16758 10044 16764 10056
rect 16715 10016 16764 10044
rect 16715 10013 16727 10016
rect 16669 10007 16727 10013
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10013 17187 10047
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 17129 10007 17187 10013
rect 11422 9976 11428 9988
rect 10888 9948 11428 9976
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 11606 9936 11612 9988
rect 11664 9936 11670 9988
rect 12897 9979 12955 9985
rect 12897 9945 12909 9979
rect 12943 9945 12955 9979
rect 16592 9976 16620 10004
rect 17144 9976 17172 10007
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 19058 10004 19064 10056
rect 19116 10044 19122 10056
rect 19392 10047 19450 10053
rect 19392 10044 19404 10047
rect 19116 10016 19404 10044
rect 19116 10004 19122 10016
rect 19392 10013 19404 10016
rect 19438 10013 19450 10047
rect 19392 10007 19450 10013
rect 21910 10004 21916 10056
rect 21968 10044 21974 10056
rect 22005 10047 22063 10053
rect 22005 10044 22017 10047
rect 21968 10016 22017 10044
rect 21968 10004 21974 10016
rect 22005 10013 22017 10016
rect 22051 10013 22063 10047
rect 22005 10007 22063 10013
rect 18230 9976 18236 9988
rect 16592 9948 17172 9976
rect 18143 9948 18236 9976
rect 12897 9939 12955 9945
rect 10594 9868 10600 9920
rect 10652 9908 10658 9920
rect 12912 9908 12940 9939
rect 18230 9936 18236 9948
rect 18288 9976 18294 9988
rect 19242 9976 19248 9988
rect 18288 9948 18920 9976
rect 19203 9948 19248 9976
rect 18288 9936 18294 9948
rect 10652 9880 12940 9908
rect 10652 9868 10658 9880
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14277 9911 14335 9917
rect 14277 9908 14289 9911
rect 14240 9880 14289 9908
rect 14240 9868 14246 9880
rect 14277 9877 14289 9880
rect 14323 9908 14335 9911
rect 17126 9908 17132 9920
rect 14323 9880 17132 9908
rect 14323 9877 14335 9880
rect 14277 9871 14335 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17402 9868 17408 9920
rect 17460 9908 17466 9920
rect 17589 9911 17647 9917
rect 17589 9908 17601 9911
rect 17460 9880 17601 9908
rect 17460 9868 17466 9880
rect 17589 9877 17601 9880
rect 17635 9877 17647 9911
rect 17589 9871 17647 9877
rect 18601 9911 18659 9917
rect 18601 9877 18613 9911
rect 18647 9908 18659 9911
rect 18782 9908 18788 9920
rect 18647 9880 18788 9908
rect 18647 9877 18659 9880
rect 18601 9871 18659 9877
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 18892 9908 18920 9948
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 19981 9979 20039 9985
rect 19981 9945 19993 9979
rect 20027 9976 20039 9979
rect 21726 9976 21732 9988
rect 20027 9948 21732 9976
rect 20027 9945 20039 9948
rect 19981 9939 20039 9945
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 22278 9976 22284 9988
rect 22239 9948 22284 9976
rect 22278 9936 22284 9948
rect 22336 9936 22342 9988
rect 24026 9976 24032 9988
rect 19334 9908 19340 9920
rect 18892 9880 19340 9908
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 22646 9868 22652 9920
rect 22704 9908 22710 9920
rect 22756 9908 22784 9976
rect 23987 9948 24032 9976
rect 24026 9936 24032 9948
rect 24084 9936 24090 9988
rect 22704 9880 22784 9908
rect 22704 9868 22710 9880
rect 1104 9818 28336 9840
rect 1104 9766 1782 9818
rect 1834 9766 1846 9818
rect 1898 9766 1910 9818
rect 1962 9766 1974 9818
rect 2026 9766 4782 9818
rect 4834 9766 4846 9818
rect 4898 9766 4910 9818
rect 4962 9766 4974 9818
rect 5026 9766 7782 9818
rect 7834 9766 7846 9818
rect 7898 9766 7910 9818
rect 7962 9766 7974 9818
rect 8026 9766 10782 9818
rect 10834 9766 10846 9818
rect 10898 9766 10910 9818
rect 10962 9766 10974 9818
rect 11026 9766 13782 9818
rect 13834 9766 13846 9818
rect 13898 9766 13910 9818
rect 13962 9766 13974 9818
rect 14026 9766 16782 9818
rect 16834 9766 16846 9818
rect 16898 9766 16910 9818
rect 16962 9766 16974 9818
rect 17026 9766 19782 9818
rect 19834 9766 19846 9818
rect 19898 9766 19910 9818
rect 19962 9766 19974 9818
rect 20026 9766 22782 9818
rect 22834 9766 22846 9818
rect 22898 9766 22910 9818
rect 22962 9766 22974 9818
rect 23026 9766 25782 9818
rect 25834 9766 25846 9818
rect 25898 9766 25910 9818
rect 25962 9766 25974 9818
rect 26026 9766 28336 9818
rect 1104 9744 28336 9766
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 7377 9707 7435 9713
rect 7377 9704 7389 9707
rect 7064 9676 7389 9704
rect 7064 9664 7070 9676
rect 7377 9673 7389 9676
rect 7423 9704 7435 9707
rect 9769 9707 9827 9713
rect 7423 9676 7788 9704
rect 7423 9673 7435 9676
rect 7377 9667 7435 9673
rect 7760 9645 7788 9676
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 9858 9704 9864 9716
rect 9815 9676 9864 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 11701 9707 11759 9713
rect 11701 9704 11713 9707
rect 11204 9676 11713 9704
rect 11204 9664 11210 9676
rect 11701 9673 11713 9676
rect 11747 9673 11759 9707
rect 13630 9704 13636 9716
rect 13591 9676 13636 9704
rect 11701 9667 11759 9673
rect 13630 9664 13636 9676
rect 13688 9704 13694 9716
rect 14090 9704 14096 9716
rect 13688 9676 14096 9704
rect 13688 9664 13694 9676
rect 14090 9664 14096 9676
rect 14148 9664 14154 9716
rect 14461 9707 14519 9713
rect 14461 9673 14473 9707
rect 14507 9704 14519 9707
rect 14550 9704 14556 9716
rect 14507 9676 14556 9704
rect 14507 9673 14519 9676
rect 14461 9667 14519 9673
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 15289 9707 15347 9713
rect 15289 9673 15301 9707
rect 15335 9704 15347 9707
rect 16206 9704 16212 9716
rect 15335 9676 16212 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 17586 9704 17592 9716
rect 17499 9676 17592 9704
rect 17586 9664 17592 9676
rect 17644 9704 17650 9716
rect 18230 9704 18236 9716
rect 17644 9676 18236 9704
rect 17644 9664 17650 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 21177 9707 21235 9713
rect 21177 9673 21189 9707
rect 21223 9673 21235 9707
rect 21177 9667 21235 9673
rect 7745 9639 7803 9645
rect 7745 9605 7757 9639
rect 7791 9605 7803 9639
rect 7745 9599 7803 9605
rect 11057 9639 11115 9645
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 11882 9636 11888 9648
rect 11103 9608 11888 9636
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 11882 9596 11888 9608
rect 11940 9596 11946 9648
rect 15654 9636 15660 9648
rect 15615 9608 15660 9636
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 18966 9596 18972 9648
rect 19024 9636 19030 9648
rect 20165 9639 20223 9645
rect 20165 9636 20177 9639
rect 19024 9608 20177 9636
rect 19024 9596 19030 9608
rect 20165 9605 20177 9608
rect 20211 9636 20223 9639
rect 20533 9639 20591 9645
rect 20533 9636 20545 9639
rect 20211 9608 20545 9636
rect 20211 9605 20223 9608
rect 20165 9599 20223 9605
rect 20533 9605 20545 9608
rect 20579 9636 20591 9639
rect 20806 9636 20812 9648
rect 20579 9608 20812 9636
rect 20579 9605 20591 9608
rect 20533 9599 20591 9605
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 21192 9636 21220 9667
rect 22278 9664 22284 9716
rect 22336 9704 22342 9716
rect 22373 9707 22431 9713
rect 22373 9704 22385 9707
rect 22336 9676 22385 9704
rect 22336 9664 22342 9676
rect 22373 9673 22385 9676
rect 22419 9673 22431 9707
rect 22373 9667 22431 9673
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 22741 9707 22799 9713
rect 22741 9704 22753 9707
rect 22704 9676 22753 9704
rect 22704 9664 22710 9676
rect 22741 9673 22753 9676
rect 22787 9673 22799 9707
rect 22741 9667 22799 9673
rect 22664 9636 22692 9664
rect 21192 9608 22692 9636
rect 8202 9568 8208 9580
rect 8163 9540 8208 9568
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 8496 9500 8524 9531
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 8628 9540 8673 9568
rect 8628 9528 8634 9540
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10502 9568 10508 9580
rect 9824 9540 10508 9568
rect 9824 9528 9830 9540
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10652 9540 10701 9568
rect 10652 9528 10658 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9568 12679 9571
rect 12894 9568 12900 9580
rect 12667 9540 12900 9568
rect 12667 9537 12679 9540
rect 12621 9531 12679 9537
rect 12894 9528 12900 9540
rect 12952 9528 12958 9580
rect 14458 9568 14464 9580
rect 14419 9540 14464 9568
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9568 16083 9571
rect 16298 9568 16304 9580
rect 16071 9540 16304 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 16298 9528 16304 9540
rect 16356 9568 16362 9580
rect 16356 9540 16528 9568
rect 16356 9528 16362 9540
rect 9030 9500 9036 9512
rect 8496 9472 8616 9500
rect 8991 9472 9036 9500
rect 6457 9435 6515 9441
rect 6457 9401 6469 9435
rect 6503 9432 6515 9435
rect 7466 9432 7472 9444
rect 6503 9404 7472 9432
rect 6503 9401 6515 9404
rect 6457 9395 6515 9401
rect 7466 9392 7472 9404
rect 7524 9392 7530 9444
rect 8588 9432 8616 9472
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9180 9472 9225 9500
rect 9180 9460 9186 9472
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 16114 9500 16120 9512
rect 11756 9472 16120 9500
rect 11756 9460 11762 9472
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 16500 9500 16528 9540
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16632 9540 16681 9568
rect 16632 9528 16638 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 19334 9568 19340 9580
rect 19295 9540 19340 9568
rect 16669 9531 16727 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19702 9568 19708 9580
rect 19444 9540 19708 9568
rect 17310 9500 17316 9512
rect 16500 9472 17316 9500
rect 17310 9460 17316 9472
rect 17368 9500 17374 9512
rect 19444 9500 19472 9540
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 20070 9568 20076 9580
rect 19843 9540 20076 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 17368 9472 19472 9500
rect 17368 9460 17374 9472
rect 19518 9460 19524 9512
rect 19576 9500 19582 9512
rect 19812 9500 19840 9531
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 20990 9568 20996 9580
rect 20903 9540 20996 9568
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 22646 9568 22652 9580
rect 21140 9540 22652 9568
rect 21140 9528 21146 9540
rect 22646 9528 22652 9540
rect 22704 9568 22710 9580
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22704 9540 23121 9568
rect 22704 9528 22710 9540
rect 23109 9537 23121 9540
rect 23155 9568 23167 9571
rect 24026 9568 24032 9580
rect 23155 9540 24032 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 19576 9472 19840 9500
rect 21008 9500 21036 9528
rect 21008 9472 21588 9500
rect 19576 9460 19582 9472
rect 8754 9432 8760 9444
rect 8588 9404 8760 9432
rect 8754 9392 8760 9404
rect 8812 9432 8818 9444
rect 11422 9432 11428 9444
rect 8812 9404 9996 9432
rect 11335 9404 11428 9432
rect 8812 9392 8818 9404
rect 9968 9376 9996 9404
rect 11422 9392 11428 9404
rect 11480 9432 11486 9444
rect 11882 9432 11888 9444
rect 11480 9404 11888 9432
rect 11480 9392 11486 9404
rect 11882 9392 11888 9404
rect 11940 9432 11946 9444
rect 13538 9432 13544 9444
rect 11940 9404 13544 9432
rect 11940 9392 11946 9404
rect 13538 9392 13544 9404
rect 13596 9432 13602 9444
rect 14182 9432 14188 9444
rect 13596 9404 14188 9432
rect 13596 9392 13602 9404
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 16298 9392 16304 9444
rect 16356 9432 16362 9444
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 16356 9404 16865 9432
rect 16356 9392 16362 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16853 9395 16911 9401
rect 19153 9435 19211 9441
rect 19153 9401 19165 9435
rect 19199 9432 19211 9435
rect 21174 9432 21180 9444
rect 19199 9404 21180 9432
rect 19199 9401 19211 9404
rect 19153 9395 19211 9401
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 21560 9441 21588 9472
rect 21545 9435 21603 9441
rect 21545 9401 21557 9435
rect 21591 9432 21603 9435
rect 22186 9432 22192 9444
rect 21591 9404 22192 9432
rect 21591 9401 21603 9404
rect 21545 9395 21603 9401
rect 22186 9392 22192 9404
rect 22244 9392 22250 9444
rect 7098 9364 7104 9376
rect 7059 9336 7104 9364
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 10008 9336 10057 9364
rect 10008 9324 10014 9336
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 10045 9327 10103 9333
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12805 9367 12863 9373
rect 12805 9364 12817 9367
rect 11664 9336 12817 9364
rect 11664 9324 11670 9336
rect 12805 9333 12817 9336
rect 12851 9333 12863 9367
rect 12805 9327 12863 9333
rect 16393 9367 16451 9373
rect 16393 9333 16405 9367
rect 16439 9364 16451 9367
rect 16666 9364 16672 9376
rect 16439 9336 16672 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16666 9324 16672 9336
rect 16724 9364 16730 9376
rect 17129 9367 17187 9373
rect 17129 9364 17141 9367
rect 16724 9336 17141 9364
rect 16724 9324 16730 9336
rect 17129 9333 17141 9336
rect 17175 9333 17187 9367
rect 17129 9327 17187 9333
rect 18601 9367 18659 9373
rect 18601 9333 18613 9367
rect 18647 9364 18659 9367
rect 19058 9364 19064 9376
rect 18647 9336 19064 9364
rect 18647 9333 18659 9336
rect 18601 9327 18659 9333
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 21910 9324 21916 9376
rect 21968 9364 21974 9376
rect 22005 9367 22063 9373
rect 22005 9364 22017 9367
rect 21968 9336 22017 9364
rect 21968 9324 21974 9336
rect 22005 9333 22017 9336
rect 22051 9333 22063 9367
rect 22005 9327 22063 9333
rect 1104 9274 28336 9296
rect 1104 9222 3282 9274
rect 3334 9222 3346 9274
rect 3398 9222 3410 9274
rect 3462 9222 3474 9274
rect 3526 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 6410 9274
rect 6462 9222 6474 9274
rect 6526 9222 9282 9274
rect 9334 9222 9346 9274
rect 9398 9222 9410 9274
rect 9462 9222 9474 9274
rect 9526 9222 12282 9274
rect 12334 9222 12346 9274
rect 12398 9222 12410 9274
rect 12462 9222 12474 9274
rect 12526 9222 15282 9274
rect 15334 9222 15346 9274
rect 15398 9222 15410 9274
rect 15462 9222 15474 9274
rect 15526 9222 18282 9274
rect 18334 9222 18346 9274
rect 18398 9222 18410 9274
rect 18462 9222 18474 9274
rect 18526 9222 21282 9274
rect 21334 9222 21346 9274
rect 21398 9222 21410 9274
rect 21462 9222 21474 9274
rect 21526 9222 24282 9274
rect 24334 9222 24346 9274
rect 24398 9222 24410 9274
rect 24462 9222 24474 9274
rect 24526 9222 27282 9274
rect 27334 9222 27346 9274
rect 27398 9222 27410 9274
rect 27462 9222 27474 9274
rect 27526 9222 28336 9274
rect 1104 9200 28336 9222
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7466 9160 7472 9172
rect 7423 9132 7472 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8352 9132 8493 9160
rect 8352 9120 8358 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 9030 9160 9036 9172
rect 8991 9132 9036 9160
rect 8481 9123 8539 9129
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 10965 9163 11023 9169
rect 10965 9129 10977 9163
rect 11011 9160 11023 9163
rect 11606 9160 11612 9172
rect 11011 9132 11612 9160
rect 11011 9129 11023 9132
rect 10965 9123 11023 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 13817 9163 13875 9169
rect 13817 9129 13829 9163
rect 13863 9160 13875 9163
rect 14274 9160 14280 9172
rect 13863 9132 14280 9160
rect 13863 9129 13875 9132
rect 13817 9123 13875 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14458 9160 14464 9172
rect 14419 9132 14464 9160
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 16264 9132 16313 9160
rect 16264 9120 16270 9132
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 16301 9123 16359 9129
rect 19521 9163 19579 9169
rect 19521 9129 19533 9163
rect 19567 9160 19579 9163
rect 19610 9160 19616 9172
rect 19567 9132 19616 9160
rect 19567 9129 19579 9132
rect 19521 9123 19579 9129
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 19702 9120 19708 9172
rect 19760 9160 19766 9172
rect 20165 9163 20223 9169
rect 20165 9160 20177 9163
rect 19760 9132 20177 9160
rect 19760 9120 19766 9132
rect 20165 9129 20177 9132
rect 20211 9129 20223 9163
rect 22278 9160 22284 9172
rect 22239 9132 22284 9160
rect 20165 9123 20223 9129
rect 22278 9120 22284 9132
rect 22336 9120 22342 9172
rect 6917 9095 6975 9101
rect 6917 9061 6929 9095
rect 6963 9092 6975 9095
rect 8202 9092 8208 9104
rect 6963 9064 8208 9092
rect 6963 9061 6975 9064
rect 6917 9055 6975 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 11241 9095 11299 9101
rect 11241 9092 11253 9095
rect 10560 9064 11253 9092
rect 10560 9052 10566 9064
rect 11241 9061 11253 9064
rect 11287 9061 11299 9095
rect 11241 9055 11299 9061
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 9024 6607 9027
rect 9122 9024 9128 9036
rect 6595 8996 9128 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 10410 9024 10416 9036
rect 10371 8996 10416 9024
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 16022 8984 16028 9036
rect 16080 9024 16086 9036
rect 16482 9024 16488 9036
rect 16080 8996 16488 9024
rect 16080 8984 16086 8996
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 17402 9024 17408 9036
rect 17363 8996 17408 9024
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 19150 9024 19156 9036
rect 19111 8996 19156 9024
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 21082 9024 21088 9036
rect 21043 8996 21088 9024
rect 21082 8984 21088 8996
rect 21140 8984 21146 9036
rect 7190 8956 7196 8968
rect 7151 8928 7196 8956
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 8202 8956 8208 8968
rect 8163 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 10045 8959 10103 8965
rect 8352 8928 8397 8956
rect 8352 8916 8358 8928
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10318 8956 10324 8968
rect 10091 8928 10324 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11940 8928 12081 8956
rect 11940 8916 11946 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8956 13691 8959
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13679 8928 14105 8956
rect 13679 8925 13691 8928
rect 13633 8919 13691 8925
rect 14093 8925 14105 8928
rect 14139 8956 14151 8959
rect 14366 8956 14372 8968
rect 14139 8928 14372 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 15102 8916 15108 8968
rect 15160 8956 15166 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15160 8928 15485 8956
rect 15160 8916 15166 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15562 8916 15568 8968
rect 15620 8956 15626 8968
rect 17126 8956 17132 8968
rect 15620 8928 15665 8956
rect 17087 8928 17132 8956
rect 15620 8916 15626 8928
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 21174 8916 21180 8968
rect 21232 8956 21238 8968
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 21232 8928 21281 8956
rect 21232 8916 21238 8928
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 21818 8916 21824 8968
rect 21876 8956 21882 8968
rect 22002 8956 22008 8968
rect 21876 8928 21921 8956
rect 21963 8928 22008 8956
rect 21876 8916 21882 8928
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 7837 8891 7895 8897
rect 7837 8857 7849 8891
rect 7883 8888 7895 8891
rect 8570 8888 8576 8900
rect 7883 8860 8576 8888
rect 7883 8857 7895 8860
rect 7837 8851 7895 8857
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 9858 8888 9864 8900
rect 9819 8860 9864 8888
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 12710 8888 12716 8900
rect 12671 8860 12716 8888
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 16022 8888 16028 8900
rect 15983 8860 16028 8888
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 17862 8848 17868 8900
rect 17920 8848 17926 8900
rect 6178 8820 6184 8832
rect 6139 8792 6184 8820
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12952 8792 13001 8820
rect 12952 8780 12958 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 14918 8820 14924 8832
rect 14879 8792 14924 8820
rect 12989 8783 13047 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16632 8792 16681 8820
rect 16632 8780 16638 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 19889 8823 19947 8829
rect 19889 8789 19901 8823
rect 19935 8820 19947 8823
rect 20254 8820 20260 8832
rect 19935 8792 20260 8820
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 1104 8730 28336 8752
rect 1104 8678 1782 8730
rect 1834 8678 1846 8730
rect 1898 8678 1910 8730
rect 1962 8678 1974 8730
rect 2026 8678 4782 8730
rect 4834 8678 4846 8730
rect 4898 8678 4910 8730
rect 4962 8678 4974 8730
rect 5026 8678 7782 8730
rect 7834 8678 7846 8730
rect 7898 8678 7910 8730
rect 7962 8678 7974 8730
rect 8026 8678 10782 8730
rect 10834 8678 10846 8730
rect 10898 8678 10910 8730
rect 10962 8678 10974 8730
rect 11026 8678 13782 8730
rect 13834 8678 13846 8730
rect 13898 8678 13910 8730
rect 13962 8678 13974 8730
rect 14026 8678 16782 8730
rect 16834 8678 16846 8730
rect 16898 8678 16910 8730
rect 16962 8678 16974 8730
rect 17026 8678 19782 8730
rect 19834 8678 19846 8730
rect 19898 8678 19910 8730
rect 19962 8678 19974 8730
rect 20026 8678 22782 8730
rect 22834 8678 22846 8730
rect 22898 8678 22910 8730
rect 22962 8678 22974 8730
rect 23026 8678 25782 8730
rect 25834 8678 25846 8730
rect 25898 8678 25910 8730
rect 25962 8678 25974 8730
rect 26026 8678 28336 8730
rect 1104 8656 28336 8678
rect 8202 8616 8208 8628
rect 8163 8588 8208 8616
rect 8202 8576 8208 8588
rect 8260 8616 8266 8628
rect 15562 8616 15568 8628
rect 8260 8588 10088 8616
rect 8260 8576 8266 8588
rect 9030 8508 9036 8560
rect 9088 8548 9094 8560
rect 9125 8551 9183 8557
rect 9125 8548 9137 8551
rect 9088 8520 9137 8548
rect 9088 8508 9094 8520
rect 9125 8517 9137 8520
rect 9171 8517 9183 8551
rect 9125 8511 9183 8517
rect 10060 8492 10088 8588
rect 10704 8588 15568 8616
rect 10704 8557 10732 8588
rect 15562 8576 15568 8588
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 17184 8588 17417 8616
rect 17184 8576 17190 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 21729 8619 21787 8625
rect 21729 8616 21741 8619
rect 21232 8588 21741 8616
rect 21232 8576 21238 8588
rect 21729 8585 21741 8588
rect 21775 8585 21787 8619
rect 21729 8579 21787 8585
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22097 8619 22155 8625
rect 22097 8616 22109 8619
rect 22060 8588 22109 8616
rect 22060 8576 22066 8588
rect 22097 8585 22109 8588
rect 22143 8585 22155 8619
rect 22097 8579 22155 8585
rect 22646 8576 22652 8628
rect 22704 8616 22710 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22704 8588 22845 8616
rect 22704 8576 22710 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 10689 8551 10747 8557
rect 10689 8517 10701 8551
rect 10735 8517 10747 8551
rect 10689 8511 10747 8517
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 12952 8520 13768 8548
rect 12952 8508 12958 8520
rect 14918 8508 14924 8560
rect 14976 8548 14982 8560
rect 14976 8520 18460 8548
rect 14976 8508 14982 8520
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8449 8631 8483
rect 8573 8443 8631 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 8938 8480 8944 8492
rect 8803 8452 8944 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 8588 8412 8616 8443
rect 8938 8440 8944 8452
rect 8996 8480 9002 8492
rect 9950 8480 9956 8492
rect 8996 8452 9812 8480
rect 9911 8452 9956 8480
rect 8996 8440 9002 8452
rect 9784 8412 9812 8452
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10229 8483 10287 8489
rect 10100 8452 10193 8480
rect 10100 8440 10106 8452
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10594 8480 10600 8492
rect 10275 8452 10600 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10244 8412 10272 8443
rect 10594 8440 10600 8452
rect 10652 8480 10658 8492
rect 10965 8483 11023 8489
rect 10965 8480 10977 8483
rect 10652 8452 10977 8480
rect 10652 8440 10658 8452
rect 10965 8449 10977 8452
rect 11011 8480 11023 8483
rect 11698 8480 11704 8492
rect 11011 8452 11704 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12768 8452 13001 8480
rect 12768 8440 12774 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 16298 8480 16304 8492
rect 15160 8452 16304 8480
rect 15160 8440 15166 8452
rect 16298 8440 16304 8452
rect 16356 8480 16362 8492
rect 16485 8483 16543 8489
rect 16485 8480 16497 8483
rect 16356 8452 16497 8480
rect 16356 8440 16362 8452
rect 16485 8449 16497 8452
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 18138 8480 18144 8492
rect 17175 8452 18144 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 18138 8440 18144 8452
rect 18196 8480 18202 8492
rect 18432 8489 18460 8520
rect 20806 8508 20812 8560
rect 20864 8548 20870 8560
rect 21361 8551 21419 8557
rect 21361 8548 21373 8551
rect 20864 8520 21373 8548
rect 20864 8508 20870 8520
rect 21361 8517 21373 8520
rect 21407 8548 21419 8551
rect 21634 8548 21640 8560
rect 21407 8520 21640 8548
rect 21407 8517 21419 8520
rect 21361 8511 21419 8517
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18196 8452 18245 8480
rect 18196 8440 18202 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8480 18475 8483
rect 19150 8480 19156 8492
rect 18463 8452 19156 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19610 8480 19616 8492
rect 19571 8452 19616 8480
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 19886 8480 19892 8492
rect 19847 8452 19892 8480
rect 19705 8443 19763 8449
rect 13262 8412 13268 8424
rect 8588 8384 9720 8412
rect 9784 8384 10272 8412
rect 13223 8384 13268 8412
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 7190 8276 7196 8288
rect 5776 8248 7196 8276
rect 5776 8236 5782 8248
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7926 8276 7932 8288
rect 7887 8248 7932 8276
rect 7926 8236 7932 8248
rect 7984 8276 7990 8288
rect 8294 8276 8300 8288
rect 7984 8248 8300 8276
rect 7984 8236 7990 8248
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 9692 8285 9720 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 14458 8372 14464 8424
rect 14516 8412 14522 8424
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 14516 8384 15025 8412
rect 14516 8372 14522 8384
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 19720 8412 19748 8443
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 20254 8480 20260 8492
rect 20215 8452 20260 8480
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20438 8480 20444 8492
rect 20496 8489 20502 8492
rect 20408 8452 20444 8480
rect 20438 8440 20444 8452
rect 20496 8480 20508 8489
rect 21542 8480 21548 8492
rect 20496 8452 21548 8480
rect 20496 8443 20508 8452
rect 20496 8440 20502 8443
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 15013 8375 15071 8381
rect 19168 8384 19748 8412
rect 9677 8279 9735 8285
rect 9677 8245 9689 8279
rect 9723 8276 9735 8279
rect 9858 8276 9864 8288
rect 9723 8248 9864 8276
rect 9723 8245 9735 8248
rect 9677 8239 9735 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 11882 8236 11888 8288
rect 11940 8276 11946 8288
rect 11977 8279 12035 8285
rect 11977 8276 11989 8279
rect 11940 8248 11989 8276
rect 11940 8236 11946 8248
rect 11977 8245 11989 8248
rect 12023 8245 12035 8279
rect 11977 8239 12035 8245
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 13998 8276 14004 8288
rect 12759 8248 14004 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 13998 8236 14004 8248
rect 14056 8276 14062 8288
rect 14476 8276 14504 8372
rect 14056 8248 14504 8276
rect 14056 8236 14062 8248
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15289 8279 15347 8285
rect 15289 8276 15301 8279
rect 15160 8248 15301 8276
rect 15160 8236 15166 8248
rect 15289 8245 15301 8248
rect 15335 8245 15347 8279
rect 15289 8239 15347 8245
rect 16117 8279 16175 8285
rect 16117 8245 16129 8279
rect 16163 8276 16175 8279
rect 16298 8276 16304 8288
rect 16163 8248 16304 8276
rect 16163 8245 16175 8248
rect 16117 8239 16175 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 17494 8236 17500 8288
rect 17552 8276 17558 8288
rect 18509 8279 18567 8285
rect 18509 8276 18521 8279
rect 17552 8248 18521 8276
rect 17552 8236 17558 8248
rect 18509 8245 18521 8248
rect 18555 8245 18567 8279
rect 18509 8239 18567 8245
rect 19058 8236 19064 8288
rect 19116 8276 19122 8288
rect 19168 8285 19196 8384
rect 20070 8372 20076 8424
rect 20128 8412 20134 8424
rect 20809 8415 20867 8421
rect 20809 8412 20821 8415
rect 20128 8384 20821 8412
rect 20128 8372 20134 8384
rect 20809 8381 20821 8384
rect 20855 8381 20867 8415
rect 20809 8375 20867 8381
rect 19153 8279 19211 8285
rect 19153 8276 19165 8279
rect 19116 8248 19165 8276
rect 19116 8236 19122 8248
rect 19153 8245 19165 8248
rect 19199 8245 19211 8279
rect 22462 8276 22468 8288
rect 22423 8248 22468 8276
rect 19153 8239 19211 8245
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 1104 8186 28336 8208
rect 1104 8134 3282 8186
rect 3334 8134 3346 8186
rect 3398 8134 3410 8186
rect 3462 8134 3474 8186
rect 3526 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 6410 8186
rect 6462 8134 6474 8186
rect 6526 8134 9282 8186
rect 9334 8134 9346 8186
rect 9398 8134 9410 8186
rect 9462 8134 9474 8186
rect 9526 8134 12282 8186
rect 12334 8134 12346 8186
rect 12398 8134 12410 8186
rect 12462 8134 12474 8186
rect 12526 8134 15282 8186
rect 15334 8134 15346 8186
rect 15398 8134 15410 8186
rect 15462 8134 15474 8186
rect 15526 8134 18282 8186
rect 18334 8134 18346 8186
rect 18398 8134 18410 8186
rect 18462 8134 18474 8186
rect 18526 8134 21282 8186
rect 21334 8134 21346 8186
rect 21398 8134 21410 8186
rect 21462 8134 21474 8186
rect 21526 8134 24282 8186
rect 24334 8134 24346 8186
rect 24398 8134 24410 8186
rect 24462 8134 24474 8186
rect 24526 8134 27282 8186
rect 27334 8134 27346 8186
rect 27398 8134 27410 8186
rect 27462 8134 27474 8186
rect 27526 8134 28336 8186
rect 1104 8112 28336 8134
rect 7469 8075 7527 8081
rect 7469 8041 7481 8075
rect 7515 8072 7527 8075
rect 8938 8072 8944 8084
rect 7515 8044 8944 8072
rect 7515 8041 7527 8044
rect 7469 8035 7527 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10042 8072 10048 8084
rect 10003 8044 10048 8072
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12253 8075 12311 8081
rect 12253 8041 12265 8075
rect 12299 8072 12311 8075
rect 12710 8072 12716 8084
rect 12299 8044 12716 8072
rect 12299 8041 12311 8044
rect 12253 8035 12311 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 14918 8072 14924 8084
rect 14879 8044 14924 8072
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17460 8044 17509 8072
rect 17460 8032 17466 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 18196 8044 18245 8072
rect 18196 8032 18202 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 18233 8035 18291 8041
rect 18858 8075 18916 8081
rect 18858 8041 18870 8075
rect 18904 8072 18916 8075
rect 19058 8072 19064 8084
rect 18904 8044 19064 8072
rect 18904 8041 18916 8044
rect 18858 8035 18916 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19337 8075 19395 8081
rect 19337 8041 19349 8075
rect 19383 8072 19395 8075
rect 19518 8072 19524 8084
rect 19383 8044 19524 8072
rect 19383 8041 19395 8044
rect 19337 8035 19395 8041
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 19610 8032 19616 8084
rect 19668 8072 19674 8084
rect 20441 8075 20499 8081
rect 20441 8072 20453 8075
rect 19668 8044 20453 8072
rect 19668 8032 19674 8044
rect 20441 8041 20453 8044
rect 20487 8041 20499 8075
rect 20441 8035 20499 8041
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 21818 8072 21824 8084
rect 21407 8044 21824 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21818 8032 21824 8044
rect 21876 8072 21882 8084
rect 22462 8072 22468 8084
rect 21876 8044 22468 8072
rect 21876 8032 21882 8044
rect 22462 8032 22468 8044
rect 22520 8032 22526 8084
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 12529 8007 12587 8013
rect 12529 8004 12541 8007
rect 7248 7976 12541 8004
rect 7248 7964 7254 7976
rect 12529 7973 12541 7976
rect 12575 8004 12587 8007
rect 12894 8004 12900 8016
rect 12575 7976 12900 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 18966 8004 18972 8016
rect 18927 7976 18972 8004
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 20254 7964 20260 8016
rect 20312 8004 20318 8016
rect 20312 7976 22232 8004
rect 20312 7964 20318 7976
rect 6178 7896 6184 7948
rect 6236 7936 6242 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 6236 7908 7113 7936
rect 6236 7896 6242 7908
rect 7101 7905 7113 7908
rect 7147 7936 7159 7939
rect 9950 7936 9956 7948
rect 7147 7908 9956 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 8588 7877 8616 7908
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 12989 7939 13047 7945
rect 12989 7905 13001 7939
rect 13035 7936 13047 7939
rect 13262 7936 13268 7948
rect 13035 7908 13268 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 15102 7936 15108 7948
rect 13924 7908 15108 7936
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7984 7840 8309 7868
rect 7984 7828 7990 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8938 7868 8944 7880
rect 8803 7840 8944 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 7466 7760 7472 7812
rect 7524 7800 7530 7812
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 7524 7772 7757 7800
rect 7524 7760 7530 7772
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 8312 7800 8340 7831
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 8662 7800 8668 7812
rect 8312 7772 8668 7800
rect 7745 7763 7803 7769
rect 8662 7760 8668 7772
rect 8720 7800 8726 7812
rect 10689 7803 10747 7809
rect 10689 7800 10701 7803
rect 8720 7772 10701 7800
rect 8720 7760 8726 7772
rect 10689 7769 10701 7772
rect 10735 7769 10747 7803
rect 10689 7763 10747 7769
rect 11256 7744 11284 7831
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 13924 7868 13952 7908
rect 15102 7896 15108 7908
rect 15160 7936 15166 7948
rect 15473 7939 15531 7945
rect 15473 7936 15485 7939
rect 15160 7908 15485 7936
rect 15160 7896 15166 7908
rect 15473 7905 15485 7908
rect 15519 7936 15531 7939
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15519 7908 15945 7936
rect 15519 7905 15531 7908
rect 15473 7899 15531 7905
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 19061 7939 19119 7945
rect 19061 7905 19073 7939
rect 19107 7936 19119 7939
rect 19610 7936 19616 7948
rect 19107 7908 19616 7936
rect 19107 7905 19119 7908
rect 19061 7899 19119 7905
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 21692 7908 22140 7936
rect 21692 7896 21698 7908
rect 13872 7840 13952 7868
rect 13872 7828 13878 7840
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14274 7868 14280 7880
rect 14235 7840 14280 7868
rect 14093 7831 14151 7837
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 15838 7828 15844 7880
rect 15896 7868 15902 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15896 7840 16037 7868
rect 15896 7828 15902 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 16206 7828 16212 7880
rect 16264 7868 16270 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 16264 7840 16497 7868
rect 16264 7828 16270 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16666 7868 16672 7880
rect 16623 7840 16672 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 16776 7840 17264 7868
rect 16776 7800 16804 7840
rect 17236 7812 17264 7840
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18196 7840 18705 7868
rect 18196 7828 18202 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7837 21603 7871
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 21545 7831 21603 7837
rect 17126 7800 17132 7812
rect 11440 7772 16804 7800
rect 17087 7772 17132 7800
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 9858 7732 9864 7744
rect 9171 7704 9864 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 11238 7732 11244 7744
rect 11151 7704 11244 7732
rect 11238 7692 11244 7704
rect 11296 7732 11302 7744
rect 11440 7732 11468 7772
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 17218 7760 17224 7812
rect 17276 7800 17282 7812
rect 19886 7800 19892 7812
rect 17276 7772 19892 7800
rect 17276 7760 17282 7772
rect 19886 7760 19892 7772
rect 19944 7800 19950 7812
rect 20073 7803 20131 7809
rect 20073 7800 20085 7803
rect 19944 7772 20085 7800
rect 19944 7760 19950 7772
rect 20073 7769 20085 7772
rect 20119 7800 20131 7803
rect 21560 7800 21588 7831
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22112 7877 22140 7908
rect 22204 7877 22232 7976
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 21818 7800 21824 7812
rect 20119 7772 21824 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 21818 7760 21824 7772
rect 21876 7760 21882 7812
rect 11296 7704 11468 7732
rect 11296 7692 11302 7704
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 17862 7732 17868 7744
rect 15804 7704 17868 7732
rect 15804 7692 15810 7704
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 19705 7735 19763 7741
rect 19705 7732 19717 7735
rect 18748 7704 19717 7732
rect 18748 7692 18754 7704
rect 19705 7701 19717 7704
rect 19751 7732 19763 7735
rect 20438 7732 20444 7744
rect 19751 7704 20444 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 1104 7642 28336 7664
rect 1104 7590 1782 7642
rect 1834 7590 1846 7642
rect 1898 7590 1910 7642
rect 1962 7590 1974 7642
rect 2026 7590 4782 7642
rect 4834 7590 4846 7642
rect 4898 7590 4910 7642
rect 4962 7590 4974 7642
rect 5026 7590 7782 7642
rect 7834 7590 7846 7642
rect 7898 7590 7910 7642
rect 7962 7590 7974 7642
rect 8026 7590 10782 7642
rect 10834 7590 10846 7642
rect 10898 7590 10910 7642
rect 10962 7590 10974 7642
rect 11026 7590 13782 7642
rect 13834 7590 13846 7642
rect 13898 7590 13910 7642
rect 13962 7590 13974 7642
rect 14026 7590 16782 7642
rect 16834 7590 16846 7642
rect 16898 7590 16910 7642
rect 16962 7590 16974 7642
rect 17026 7590 19782 7642
rect 19834 7590 19846 7642
rect 19898 7590 19910 7642
rect 19962 7590 19974 7642
rect 20026 7590 22782 7642
rect 22834 7590 22846 7642
rect 22898 7590 22910 7642
rect 22962 7590 22974 7642
rect 23026 7590 25782 7642
rect 25834 7590 25846 7642
rect 25898 7590 25910 7642
rect 25962 7590 25974 7642
rect 26026 7590 28336 7642
rect 1104 7568 28336 7590
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 8938 7528 8944 7540
rect 8899 7500 8944 7528
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 10781 7531 10839 7537
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 11238 7528 11244 7540
rect 10827 7500 11244 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13630 7528 13636 7540
rect 13587 7500 13636 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14274 7528 14280 7540
rect 14235 7500 14280 7528
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 16114 7528 16120 7540
rect 16075 7500 16120 7528
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17218 7528 17224 7540
rect 17175 7500 17224 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 18138 7488 18144 7540
rect 18196 7528 18202 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18196 7500 18337 7528
rect 18196 7488 18202 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 19610 7528 19616 7540
rect 18325 7491 18383 7497
rect 19444 7500 19616 7528
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 10100 7432 10149 7460
rect 10100 7420 10106 7432
rect 10137 7429 10149 7432
rect 10183 7429 10195 7463
rect 10137 7423 10195 7429
rect 14829 7463 14887 7469
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 15105 7463 15163 7469
rect 15105 7460 15117 7463
rect 14875 7432 15117 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 15105 7429 15117 7432
rect 15151 7460 15163 7463
rect 15838 7460 15844 7472
rect 15151 7432 15844 7460
rect 15151 7429 15163 7432
rect 15105 7423 15163 7429
rect 15838 7420 15844 7432
rect 15896 7420 15902 7472
rect 16390 7420 16396 7472
rect 16448 7460 16454 7472
rect 19444 7469 19472 7500
rect 19610 7488 19616 7500
rect 19668 7528 19674 7540
rect 19705 7531 19763 7537
rect 19705 7528 19717 7531
rect 19668 7500 19717 7528
rect 19668 7488 19674 7500
rect 19705 7497 19717 7500
rect 19751 7497 19763 7531
rect 19705 7491 19763 7497
rect 21726 7488 21732 7540
rect 21784 7528 21790 7540
rect 22741 7531 22799 7537
rect 22741 7528 22753 7531
rect 21784 7500 22753 7528
rect 21784 7488 21790 7500
rect 22741 7497 22753 7500
rect 22787 7497 22799 7531
rect 22741 7491 22799 7497
rect 17405 7463 17463 7469
rect 17405 7460 17417 7463
rect 16448 7432 17417 7460
rect 16448 7420 16454 7432
rect 17405 7429 17417 7432
rect 17451 7429 17463 7463
rect 17405 7423 17463 7429
rect 19429 7463 19487 7469
rect 19429 7429 19441 7463
rect 19475 7429 19487 7463
rect 21818 7460 21824 7472
rect 21779 7432 21824 7460
rect 19429 7423 19487 7429
rect 21818 7420 21824 7432
rect 21876 7420 21882 7472
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 7524 7364 7573 7392
rect 7524 7352 7530 7364
rect 7561 7361 7573 7364
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 9122 7392 9128 7404
rect 8343 7364 9128 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 8312 7324 8340 7355
rect 9122 7352 9128 7364
rect 9180 7392 9186 7404
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9180 7364 9505 7392
rect 9180 7352 9186 7364
rect 9493 7361 9505 7364
rect 9539 7392 9551 7395
rect 10318 7392 10324 7404
rect 9539 7364 10324 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 11756 7364 12725 7392
rect 11756 7352 11762 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 13722 7392 13728 7404
rect 12952 7364 13728 7392
rect 12952 7352 12958 7364
rect 13722 7352 13728 7364
rect 13780 7392 13786 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13780 7364 13829 7392
rect 13780 7352 13786 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 15562 7392 15568 7404
rect 15523 7364 15568 7392
rect 13817 7355 13875 7361
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17034 7392 17040 7404
rect 16991 7364 17040 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17034 7352 17040 7364
rect 17092 7392 17098 7404
rect 17494 7392 17500 7404
rect 17092 7364 17500 7392
rect 17092 7352 17098 7364
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 20990 7352 20996 7404
rect 21048 7392 21054 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 21048 7364 21281 7392
rect 21048 7352 21054 7364
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21726 7392 21732 7404
rect 21499 7364 21732 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 22278 7392 22284 7404
rect 22239 7364 22284 7392
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 7331 7296 8340 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 9950 7284 9956 7336
rect 10008 7324 10014 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10008 7296 11069 7324
rect 10008 7284 10014 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 12618 7324 12624 7336
rect 12579 7296 12624 7324
rect 11057 7287 11115 7293
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 20809 7327 20867 7333
rect 20809 7324 20821 7327
rect 20680 7296 20821 7324
rect 20680 7284 20686 7296
rect 20809 7293 20821 7296
rect 20855 7324 20867 7327
rect 21174 7324 21180 7336
rect 20855 7296 21180 7324
rect 20855 7293 20867 7296
rect 20809 7287 20867 7293
rect 21174 7284 21180 7296
rect 21232 7284 21238 7336
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 13446 7256 13452 7268
rect 11747 7228 13452 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 13446 7216 13452 7228
rect 13504 7256 13510 7268
rect 14274 7256 14280 7268
rect 13504 7228 14280 7256
rect 13504 7216 13510 7228
rect 14274 7216 14280 7228
rect 14332 7216 14338 7268
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 7653 7191 7711 7197
rect 7653 7188 7665 7191
rect 7616 7160 7665 7188
rect 7616 7148 7622 7160
rect 7653 7157 7665 7160
rect 7699 7157 7711 7191
rect 12066 7188 12072 7200
rect 12027 7160 12072 7188
rect 7653 7151 7711 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 13136 7160 14013 7188
rect 13136 7148 13142 7160
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 14001 7151 14059 7157
rect 15930 7148 15936 7200
rect 15988 7188 15994 7200
rect 16485 7191 16543 7197
rect 16485 7188 16497 7191
rect 15988 7160 16497 7188
rect 15988 7148 15994 7160
rect 16485 7157 16497 7160
rect 16531 7188 16543 7191
rect 16666 7188 16672 7200
rect 16531 7160 16672 7188
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 20530 7188 20536 7200
rect 20491 7160 20536 7188
rect 20530 7148 20536 7160
rect 20588 7148 20594 7200
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 21910 7188 21916 7200
rect 21232 7160 21916 7188
rect 21232 7148 21238 7160
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 1104 7098 28336 7120
rect 1104 7046 3282 7098
rect 3334 7046 3346 7098
rect 3398 7046 3410 7098
rect 3462 7046 3474 7098
rect 3526 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 6410 7098
rect 6462 7046 6474 7098
rect 6526 7046 9282 7098
rect 9334 7046 9346 7098
rect 9398 7046 9410 7098
rect 9462 7046 9474 7098
rect 9526 7046 12282 7098
rect 12334 7046 12346 7098
rect 12398 7046 12410 7098
rect 12462 7046 12474 7098
rect 12526 7046 15282 7098
rect 15334 7046 15346 7098
rect 15398 7046 15410 7098
rect 15462 7046 15474 7098
rect 15526 7046 18282 7098
rect 18334 7046 18346 7098
rect 18398 7046 18410 7098
rect 18462 7046 18474 7098
rect 18526 7046 21282 7098
rect 21334 7046 21346 7098
rect 21398 7046 21410 7098
rect 21462 7046 21474 7098
rect 21526 7046 24282 7098
rect 24334 7046 24346 7098
rect 24398 7046 24410 7098
rect 24462 7046 24474 7098
rect 24526 7046 27282 7098
rect 27334 7046 27346 7098
rect 27398 7046 27410 7098
rect 27462 7046 27474 7098
rect 27526 7046 28336 7098
rect 1104 7024 28336 7046
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 14182 6984 14188 6996
rect 13780 6956 14188 6984
rect 13780 6944 13786 6956
rect 14182 6944 14188 6956
rect 14240 6984 14246 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 14240 6956 14657 6984
rect 14240 6944 14246 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 17034 6984 17040 6996
rect 16995 6956 17040 6984
rect 14645 6947 14703 6953
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 17497 6987 17555 6993
rect 17497 6953 17509 6987
rect 17543 6984 17555 6987
rect 18966 6984 18972 6996
rect 17543 6956 18972 6984
rect 17543 6953 17555 6956
rect 17497 6947 17555 6953
rect 18966 6944 18972 6956
rect 19024 6944 19030 6996
rect 20254 6944 20260 6996
rect 20312 6984 20318 6996
rect 20441 6987 20499 6993
rect 20441 6984 20453 6987
rect 20312 6956 20453 6984
rect 20312 6944 20318 6956
rect 20441 6953 20453 6956
rect 20487 6953 20499 6987
rect 20441 6947 20499 6953
rect 15562 6916 15568 6928
rect 15523 6888 15568 6916
rect 15562 6876 15568 6888
rect 15620 6876 15626 6928
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 18417 6919 18475 6925
rect 18417 6916 18429 6919
rect 15896 6888 18429 6916
rect 15896 6876 15902 6888
rect 18417 6885 18429 6888
rect 18463 6916 18475 6919
rect 19058 6916 19064 6928
rect 18463 6888 19064 6916
rect 18463 6885 18475 6888
rect 18417 6879 18475 6885
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 7650 6848 7656 6860
rect 6687 6820 7656 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 7650 6808 7656 6820
rect 7708 6848 7714 6860
rect 12069 6851 12127 6857
rect 7708 6820 7972 6848
rect 7708 6808 7714 6820
rect 6730 6740 6736 6792
rect 6788 6780 6794 6792
rect 7558 6780 7564 6792
rect 6788 6752 7564 6780
rect 6788 6740 6794 6752
rect 7558 6740 7564 6752
rect 7616 6780 7622 6792
rect 7944 6789 7972 6820
rect 12069 6817 12081 6851
rect 12115 6848 12127 6851
rect 12618 6848 12624 6860
rect 12115 6820 12624 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12618 6808 12624 6820
rect 12676 6848 12682 6860
rect 13170 6848 13176 6860
rect 12676 6820 13176 6848
rect 12676 6808 12682 6820
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 14332 6820 14381 6848
rect 14332 6808 14338 6820
rect 14369 6817 14381 6820
rect 14415 6817 14427 6851
rect 14369 6811 14427 6817
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16298 6848 16304 6860
rect 16071 6820 16304 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 19150 6808 19156 6860
rect 19208 6848 19214 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 19208 6820 19257 6848
rect 19208 6808 19214 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 19705 6851 19763 6857
rect 19705 6848 19717 6851
rect 19576 6820 19717 6848
rect 19576 6808 19582 6820
rect 19705 6817 19717 6820
rect 19751 6817 19763 6851
rect 20070 6848 20076 6860
rect 19705 6811 19763 6817
rect 19812 6820 20076 6848
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7616 6752 7757 6780
rect 7616 6740 7622 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 8110 6780 8116 6792
rect 8071 6752 8116 6780
rect 7929 6743 7987 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8570 6780 8576 6792
rect 8531 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 10502 6780 10508 6792
rect 8720 6752 8765 6780
rect 10463 6752 10508 6780
rect 8720 6740 8726 6752
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 12345 6783 12403 6789
rect 12345 6780 12357 6783
rect 11940 6752 12357 6780
rect 11940 6740 11946 6752
rect 12345 6749 12357 6752
rect 12391 6749 12403 6783
rect 12345 6743 12403 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6780 17831 6783
rect 18138 6780 18144 6792
rect 17819 6752 18144 6780
rect 17819 6749 17831 6752
rect 17773 6743 17831 6749
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 7374 6712 7380 6724
rect 7331 6684 7380 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 9858 6672 9864 6724
rect 9916 6712 9922 6724
rect 10045 6715 10103 6721
rect 10045 6712 10057 6715
rect 9916 6684 10057 6712
rect 9916 6672 9922 6684
rect 10045 6681 10057 6684
rect 10091 6681 10103 6715
rect 12618 6712 12624 6724
rect 12579 6684 12624 6712
rect 10045 6675 10103 6681
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 13078 6672 13084 6724
rect 13136 6672 13142 6724
rect 15930 6672 15936 6724
rect 15988 6712 15994 6724
rect 16132 6712 16160 6743
rect 18138 6740 18144 6752
rect 18196 6780 18202 6792
rect 18598 6780 18604 6792
rect 18196 6752 18604 6780
rect 18196 6740 18202 6752
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19812 6789 19840 6820
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 21082 6848 21088 6860
rect 20588 6820 21088 6848
rect 20588 6808 20594 6820
rect 21082 6808 21088 6820
rect 21140 6848 21146 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21140 6820 21465 6848
rect 21140 6808 21146 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 21818 6808 21824 6860
rect 21876 6848 21882 6860
rect 23201 6851 23259 6857
rect 23201 6848 23213 6851
rect 21876 6820 23213 6848
rect 21876 6808 21882 6820
rect 23201 6817 23213 6820
rect 23247 6848 23259 6851
rect 23477 6851 23535 6857
rect 23477 6848 23489 6851
rect 23247 6820 23489 6848
rect 23247 6817 23259 6820
rect 23201 6811 23259 6817
rect 23477 6817 23489 6820
rect 23523 6817 23535 6851
rect 23477 6811 23535 6817
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19392 6752 19441 6780
rect 19392 6740 19398 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 21174 6780 21180 6792
rect 21135 6752 21180 6780
rect 19797 6743 19855 6749
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 15988 6684 16160 6712
rect 15988 6672 15994 6684
rect 17586 6672 17592 6724
rect 17644 6712 17650 6724
rect 21542 6712 21548 6724
rect 17644 6684 21548 6712
rect 17644 6672 17650 6684
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 22462 6672 22468 6724
rect 22520 6672 22526 6724
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6644 7067 6647
rect 7558 6644 7564 6656
rect 7055 6616 7564 6644
rect 7055 6613 7067 6616
rect 7009 6607 7067 6613
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9217 6647 9275 6653
rect 9217 6644 9229 6647
rect 9180 6616 9229 6644
rect 9180 6604 9186 6616
rect 9217 6613 9229 6616
rect 9263 6613 9275 6647
rect 11146 6644 11152 6656
rect 11107 6616 11152 6644
rect 9217 6607 9275 6613
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11698 6644 11704 6656
rect 11659 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 17957 6647 18015 6653
rect 17957 6644 17969 6647
rect 16540 6616 17969 6644
rect 16540 6604 16546 6616
rect 17957 6613 17969 6616
rect 18003 6644 18015 6647
rect 18874 6644 18880 6656
rect 18003 6616 18880 6644
rect 18003 6613 18015 6616
rect 17957 6607 18015 6613
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 1104 6554 28336 6576
rect 1104 6502 1782 6554
rect 1834 6502 1846 6554
rect 1898 6502 1910 6554
rect 1962 6502 1974 6554
rect 2026 6502 4782 6554
rect 4834 6502 4846 6554
rect 4898 6502 4910 6554
rect 4962 6502 4974 6554
rect 5026 6502 7782 6554
rect 7834 6502 7846 6554
rect 7898 6502 7910 6554
rect 7962 6502 7974 6554
rect 8026 6502 10782 6554
rect 10834 6502 10846 6554
rect 10898 6502 10910 6554
rect 10962 6502 10974 6554
rect 11026 6502 13782 6554
rect 13834 6502 13846 6554
rect 13898 6502 13910 6554
rect 13962 6502 13974 6554
rect 14026 6502 16782 6554
rect 16834 6502 16846 6554
rect 16898 6502 16910 6554
rect 16962 6502 16974 6554
rect 17026 6502 19782 6554
rect 19834 6502 19846 6554
rect 19898 6502 19910 6554
rect 19962 6502 19974 6554
rect 20026 6502 22782 6554
rect 22834 6502 22846 6554
rect 22898 6502 22910 6554
rect 22962 6502 22974 6554
rect 23026 6502 25782 6554
rect 25834 6502 25846 6554
rect 25898 6502 25910 6554
rect 25962 6502 25974 6554
rect 26026 6502 28336 6554
rect 1104 6480 28336 6502
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 7190 6440 7196 6452
rect 5951 6412 7196 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 7190 6400 7196 6412
rect 7248 6440 7254 6452
rect 9674 6440 9680 6452
rect 7248 6412 7880 6440
rect 9587 6412 9680 6440
rect 7248 6400 7254 6412
rect 7852 6344 7880 6412
rect 9674 6400 9680 6412
rect 9732 6440 9738 6452
rect 10502 6440 10508 6452
rect 9732 6412 10508 6440
rect 9732 6400 9738 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6440 11759 6443
rect 13078 6440 13084 6452
rect 11747 6412 13084 6440
rect 11747 6409 11759 6412
rect 11701 6403 11759 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 14829 6443 14887 6449
rect 14829 6409 14841 6443
rect 14875 6440 14887 6443
rect 17586 6440 17592 6452
rect 14875 6412 17592 6440
rect 14875 6409 14887 6412
rect 14829 6403 14887 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 20070 6440 20076 6452
rect 17727 6412 20076 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 20070 6400 20076 6412
rect 20128 6400 20134 6452
rect 21542 6400 21548 6452
rect 21600 6440 21606 6452
rect 22278 6440 22284 6452
rect 21600 6412 22284 6440
rect 21600 6400 21606 6412
rect 22278 6400 22284 6412
rect 22336 6440 22342 6452
rect 22649 6443 22707 6449
rect 22649 6440 22661 6443
rect 22336 6412 22661 6440
rect 22336 6400 22342 6412
rect 22649 6409 22661 6412
rect 22695 6409 22707 6443
rect 22649 6403 22707 6409
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 8720 6276 9965 6304
rect 8720 6264 8726 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 10520 6304 10548 6400
rect 11330 6372 11336 6384
rect 11243 6344 11336 6372
rect 11330 6332 11336 6344
rect 11388 6372 11394 6384
rect 12894 6372 12900 6384
rect 11388 6344 12900 6372
rect 11388 6332 11394 6344
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 16316 6344 17141 6372
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10520 6276 10793 6304
rect 9953 6267 10011 6273
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 10781 6267 10839 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13446 6304 13452 6316
rect 13407 6276 13452 6304
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14424 6276 14657 6304
rect 14424 6264 14430 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 16316 6313 16344 6344
rect 17129 6341 17141 6344
rect 17175 6372 17187 6375
rect 17402 6372 17408 6384
rect 17175 6344 17408 6372
rect 17175 6341 17187 6344
rect 17129 6335 17187 6341
rect 17402 6332 17408 6344
rect 17460 6332 17466 6384
rect 19058 6372 19064 6384
rect 19019 6344 19064 6372
rect 19058 6332 19064 6344
rect 19116 6332 19122 6384
rect 19794 6332 19800 6384
rect 19852 6332 19858 6384
rect 21634 6372 21640 6384
rect 21595 6344 21640 6372
rect 21634 6332 21640 6344
rect 21692 6332 21698 6384
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 16080 6276 16313 6304
rect 16080 6264 16086 6276
rect 16301 6273 16313 6276
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16540 6276 16681 6304
rect 16540 6264 16546 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 21726 6304 21732 6316
rect 21687 6276 21732 6304
rect 16669 6267 16727 6273
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 7098 6236 7104 6248
rect 7059 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 9122 6236 9128 6248
rect 9083 6208 9128 6236
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 10502 6236 10508 6248
rect 10463 6208 10508 6236
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10965 6239 11023 6245
rect 10965 6205 10977 6239
rect 11011 6236 11023 6239
rect 11146 6236 11152 6248
rect 11011 6208 11152 6236
rect 11011 6205 11023 6208
rect 10965 6199 11023 6205
rect 9140 6168 9168 6196
rect 10980 6168 11008 6199
rect 11146 6196 11152 6208
rect 11204 6196 11210 6248
rect 12618 6236 12624 6248
rect 12579 6208 12624 6236
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6236 13599 6239
rect 14274 6236 14280 6248
rect 13587 6208 14280 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 14274 6196 14280 6208
rect 14332 6196 14338 6248
rect 16390 6236 16396 6248
rect 16351 6208 16396 6236
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6205 16819 6239
rect 16761 6199 16819 6205
rect 9140 6140 11008 6168
rect 15381 6171 15439 6177
rect 15381 6137 15393 6171
rect 15427 6168 15439 6171
rect 15930 6168 15936 6180
rect 15427 6140 15936 6168
rect 15427 6137 15439 6140
rect 15381 6131 15439 6137
rect 15930 6128 15936 6140
rect 15988 6168 15994 6180
rect 16776 6168 16804 6199
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 18656 6208 18797 6236
rect 18656 6196 18662 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 15988 6140 16804 6168
rect 15988 6128 15994 6140
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 8110 6100 8116 6112
rect 6503 6072 8116 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 11977 6103 12035 6109
rect 11977 6100 11989 6103
rect 11940 6072 11989 6100
rect 11940 6060 11946 6072
rect 11977 6069 11989 6072
rect 12023 6069 12035 6103
rect 11977 6063 12035 6069
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13909 6103 13967 6109
rect 13909 6100 13921 6103
rect 13044 6072 13921 6100
rect 13044 6060 13050 6072
rect 13909 6069 13921 6072
rect 13955 6069 13967 6103
rect 14366 6100 14372 6112
rect 14327 6072 14372 6100
rect 13909 6063 13967 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 15749 6103 15807 6109
rect 15749 6069 15761 6103
rect 15795 6100 15807 6103
rect 16114 6100 16120 6112
rect 15795 6072 16120 6100
rect 15795 6069 15807 6072
rect 15749 6063 15807 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 18196 6072 18245 6100
rect 18196 6060 18202 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 18800 6100 18828 6199
rect 19150 6196 19156 6248
rect 19208 6236 19214 6248
rect 20809 6239 20867 6245
rect 20809 6236 20821 6239
rect 19208 6208 20821 6236
rect 19208 6196 19214 6208
rect 20809 6205 20821 6208
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 21174 6100 21180 6112
rect 18800 6072 21180 6100
rect 18233 6063 18291 6069
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 1104 6010 28336 6032
rect 1104 5958 3282 6010
rect 3334 5958 3346 6010
rect 3398 5958 3410 6010
rect 3462 5958 3474 6010
rect 3526 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 6410 6010
rect 6462 5958 6474 6010
rect 6526 5958 9282 6010
rect 9334 5958 9346 6010
rect 9398 5958 9410 6010
rect 9462 5958 9474 6010
rect 9526 5958 12282 6010
rect 12334 5958 12346 6010
rect 12398 5958 12410 6010
rect 12462 5958 12474 6010
rect 12526 5958 15282 6010
rect 15334 5958 15346 6010
rect 15398 5958 15410 6010
rect 15462 5958 15474 6010
rect 15526 5958 18282 6010
rect 18334 5958 18346 6010
rect 18398 5958 18410 6010
rect 18462 5958 18474 6010
rect 18526 5958 21282 6010
rect 21334 5958 21346 6010
rect 21398 5958 21410 6010
rect 21462 5958 21474 6010
rect 21526 5958 24282 6010
rect 24334 5958 24346 6010
rect 24398 5958 24410 6010
rect 24462 5958 24474 6010
rect 24526 5958 27282 6010
rect 27334 5958 27346 6010
rect 27398 5958 27410 6010
rect 27462 5958 27474 6010
rect 27526 5958 28336 6010
rect 1104 5936 28336 5958
rect 5718 5896 5724 5908
rect 5679 5868 5724 5896
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 6730 5896 6736 5908
rect 6503 5868 6736 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 6825 5899 6883 5905
rect 6825 5865 6837 5899
rect 6871 5896 6883 5899
rect 7374 5896 7380 5908
rect 6871 5868 7380 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7708 5868 8033 5896
rect 7708 5856 7714 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8628 5868 8677 5896
rect 8628 5856 8634 5868
rect 8665 5865 8677 5868
rect 8711 5896 8723 5899
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 8711 5868 10149 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 10137 5859 10195 5865
rect 12437 5899 12495 5905
rect 12437 5865 12449 5899
rect 12483 5896 12495 5899
rect 12618 5896 12624 5908
rect 12483 5868 12624 5896
rect 12483 5865 12495 5868
rect 12437 5859 12495 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 13136 5868 14289 5896
rect 13136 5856 13142 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 15746 5896 15752 5908
rect 15707 5868 15752 5896
rect 14277 5859 14335 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 19058 5896 19064 5908
rect 18279 5868 19064 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19794 5896 19800 5908
rect 19755 5868 19800 5896
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 20312 5868 20361 5896
rect 20312 5856 20318 5868
rect 20349 5865 20361 5868
rect 20395 5896 20407 5899
rect 20990 5896 20996 5908
rect 20395 5868 20996 5896
rect 20395 5865 20407 5868
rect 20349 5859 20407 5865
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 21082 5856 21088 5908
rect 21140 5896 21146 5908
rect 21177 5899 21235 5905
rect 21177 5896 21189 5899
rect 21140 5868 21189 5896
rect 21140 5856 21146 5868
rect 21177 5865 21189 5868
rect 21223 5865 21235 5899
rect 21177 5859 21235 5865
rect 21637 5899 21695 5905
rect 21637 5865 21649 5899
rect 21683 5896 21695 5899
rect 22462 5896 22468 5908
rect 21683 5868 22468 5896
rect 21683 5865 21695 5868
rect 21637 5859 21695 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 9309 5831 9367 5837
rect 9309 5797 9321 5831
rect 9355 5828 9367 5831
rect 9674 5828 9680 5840
rect 9355 5800 9680 5828
rect 9355 5797 9367 5800
rect 9309 5791 9367 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 14921 5831 14979 5837
rect 14921 5797 14933 5831
rect 14967 5828 14979 5831
rect 16022 5828 16028 5840
rect 14967 5800 16028 5828
rect 14967 5797 14979 5800
rect 14921 5791 14979 5797
rect 16022 5788 16028 5800
rect 16080 5788 16086 5840
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10560 5732 10793 5760
rect 10560 5720 10566 5732
rect 10781 5729 10793 5732
rect 10827 5760 10839 5763
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 10827 5732 11345 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11333 5729 11345 5732
rect 11379 5760 11391 5763
rect 11974 5760 11980 5772
rect 11379 5732 11980 5760
rect 11379 5729 11391 5732
rect 11333 5723 11391 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 13078 5760 13084 5772
rect 12115 5732 13084 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 18690 5760 18696 5772
rect 13786 5732 18696 5760
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8110 5692 8116 5704
rect 7975 5664 8116 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8110 5652 8116 5664
rect 8168 5692 8174 5704
rect 9122 5692 9128 5704
rect 8168 5664 9128 5692
rect 8168 5652 8174 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 10042 5692 10048 5704
rect 10003 5664 10048 5692
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 11514 5692 11520 5704
rect 11475 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5692 11578 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 11572 5664 12909 5692
rect 11572 5652 11578 5664
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13170 5692 13176 5704
rect 13044 5664 13089 5692
rect 13131 5664 13176 5692
rect 13044 5652 13050 5664
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13786 5692 13814 5732
rect 18690 5720 18696 5732
rect 18748 5720 18754 5772
rect 18874 5760 18880 5772
rect 18835 5732 18880 5760
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 19429 5763 19487 5769
rect 19429 5729 19441 5763
rect 19475 5760 19487 5763
rect 20898 5760 20904 5772
rect 19475 5732 20904 5760
rect 19475 5729 19487 5732
rect 19429 5723 19487 5729
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 13280 5664 13814 5692
rect 7650 5584 7656 5636
rect 7708 5624 7714 5636
rect 7745 5627 7803 5633
rect 7745 5624 7757 5627
rect 7708 5596 7757 5624
rect 7708 5584 7714 5596
rect 7745 5593 7757 5596
rect 7791 5593 7803 5627
rect 7745 5587 7803 5593
rect 9030 5584 9036 5636
rect 9088 5624 9094 5636
rect 9858 5624 9864 5636
rect 9088 5596 9864 5624
rect 9088 5584 9094 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 11609 5627 11667 5633
rect 11609 5624 11621 5627
rect 11388 5596 11621 5624
rect 11388 5584 11394 5596
rect 11609 5593 11621 5596
rect 11655 5593 11667 5627
rect 11609 5587 11667 5593
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 11790 5624 11796 5636
rect 11747 5596 11796 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 11790 5584 11796 5596
rect 11848 5624 11854 5636
rect 13280 5624 13308 5664
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 14608 5664 15577 5692
rect 14608 5652 14614 5664
rect 15565 5661 15577 5664
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 17129 5695 17187 5701
rect 17129 5692 17141 5695
rect 16724 5664 17141 5692
rect 16724 5652 16730 5664
rect 17129 5661 17141 5664
rect 17175 5661 17187 5695
rect 17402 5692 17408 5704
rect 17363 5664 17408 5692
rect 17129 5655 17187 5661
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18969 5695 19027 5701
rect 18969 5661 18981 5695
rect 19015 5692 19027 5695
rect 19150 5692 19156 5704
rect 19015 5664 19156 5692
rect 19015 5661 19027 5664
rect 18969 5655 19027 5661
rect 19150 5652 19156 5664
rect 19208 5652 19214 5704
rect 11848 5596 13308 5624
rect 13633 5627 13691 5633
rect 11848 5584 11854 5596
rect 13633 5593 13645 5627
rect 13679 5624 13691 5627
rect 15102 5624 15108 5636
rect 13679 5596 15108 5624
rect 13679 5593 13691 5596
rect 13633 5587 13691 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 16577 5627 16635 5633
rect 16577 5593 16589 5627
rect 16623 5624 16635 5627
rect 19242 5624 19248 5636
rect 16623 5596 19248 5624
rect 16623 5593 16635 5596
rect 16577 5587 16635 5593
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 7156 5528 7205 5556
rect 7156 5516 7162 5528
rect 7193 5525 7205 5528
rect 7239 5556 7251 5559
rect 8846 5556 8852 5568
rect 7239 5528 8852 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 8846 5516 8852 5528
rect 8904 5516 8910 5568
rect 14001 5559 14059 5565
rect 14001 5525 14013 5559
rect 14047 5556 14059 5559
rect 14274 5556 14280 5568
rect 14047 5528 14280 5556
rect 14047 5525 14059 5528
rect 14001 5519 14059 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 16022 5556 16028 5568
rect 15983 5528 16028 5556
rect 16022 5516 16028 5528
rect 16080 5516 16086 5568
rect 16206 5516 16212 5568
rect 16264 5556 16270 5568
rect 18509 5559 18567 5565
rect 18509 5556 18521 5559
rect 16264 5528 18521 5556
rect 16264 5516 16270 5528
rect 18509 5525 18521 5528
rect 18555 5556 18567 5559
rect 18598 5556 18604 5568
rect 18555 5528 18604 5556
rect 18555 5525 18567 5528
rect 18509 5519 18567 5525
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 21910 5556 21916 5568
rect 21871 5528 21916 5556
rect 21910 5516 21916 5528
rect 21968 5556 21974 5568
rect 22281 5559 22339 5565
rect 22281 5556 22293 5559
rect 21968 5528 22293 5556
rect 21968 5516 21974 5528
rect 22281 5525 22293 5528
rect 22327 5525 22339 5559
rect 22281 5519 22339 5525
rect 1104 5466 28336 5488
rect 1104 5414 1782 5466
rect 1834 5414 1846 5466
rect 1898 5414 1910 5466
rect 1962 5414 1974 5466
rect 2026 5414 4782 5466
rect 4834 5414 4846 5466
rect 4898 5414 4910 5466
rect 4962 5414 4974 5466
rect 5026 5414 7782 5466
rect 7834 5414 7846 5466
rect 7898 5414 7910 5466
rect 7962 5414 7974 5466
rect 8026 5414 10782 5466
rect 10834 5414 10846 5466
rect 10898 5414 10910 5466
rect 10962 5414 10974 5466
rect 11026 5414 13782 5466
rect 13834 5414 13846 5466
rect 13898 5414 13910 5466
rect 13962 5414 13974 5466
rect 14026 5414 16782 5466
rect 16834 5414 16846 5466
rect 16898 5414 16910 5466
rect 16962 5414 16974 5466
rect 17026 5414 19782 5466
rect 19834 5414 19846 5466
rect 19898 5414 19910 5466
rect 19962 5414 19974 5466
rect 20026 5414 22782 5466
rect 22834 5414 22846 5466
rect 22898 5414 22910 5466
rect 22962 5414 22974 5466
rect 23026 5414 25782 5466
rect 25834 5414 25846 5466
rect 25898 5414 25910 5466
rect 25962 5414 25974 5466
rect 26026 5414 28336 5466
rect 1104 5392 28336 5414
rect 7190 5352 7196 5364
rect 7151 5324 7196 5352
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7708 5324 7757 5352
rect 7708 5312 7714 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 7745 5315 7803 5321
rect 8205 5355 8263 5361
rect 8205 5321 8217 5355
rect 8251 5352 8263 5355
rect 8662 5352 8668 5364
rect 8251 5324 8668 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9030 5352 9036 5364
rect 8991 5324 9036 5352
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10042 5352 10048 5364
rect 9907 5324 10048 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10042 5312 10048 5324
rect 10100 5352 10106 5364
rect 10318 5352 10324 5364
rect 10100 5324 10324 5352
rect 10100 5312 10106 5324
rect 10318 5312 10324 5324
rect 10376 5352 10382 5364
rect 11790 5352 11796 5364
rect 10376 5324 11796 5352
rect 10376 5312 10382 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14737 5355 14795 5361
rect 14737 5321 14749 5355
rect 14783 5352 14795 5355
rect 16482 5352 16488 5364
rect 14783 5324 16488 5352
rect 14783 5321 14795 5324
rect 14737 5315 14795 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16666 5312 16672 5364
rect 16724 5352 16730 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 16724 5324 17417 5352
rect 16724 5312 16730 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 19242 5352 19248 5364
rect 19203 5324 19248 5352
rect 17405 5315 17463 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 20898 5352 20904 5364
rect 20859 5324 20904 5352
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 21726 5352 21732 5364
rect 21687 5324 21732 5352
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 11422 5284 11428 5296
rect 10796 5256 11428 5284
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 8996 5188 9321 5216
rect 8996 5176 9002 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 10796 5225 10824 5256
rect 11422 5244 11428 5256
rect 11480 5284 11486 5296
rect 15749 5287 15807 5293
rect 11480 5256 12112 5284
rect 11480 5244 11486 5256
rect 12084 5228 12112 5256
rect 15749 5253 15761 5287
rect 15795 5284 15807 5287
rect 16022 5284 16028 5296
rect 15795 5256 16028 5284
rect 15795 5253 15807 5256
rect 15749 5247 15807 5253
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 17586 5284 17592 5296
rect 16347 5256 17592 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 17586 5244 17592 5256
rect 17644 5284 17650 5296
rect 18138 5284 18144 5296
rect 17644 5256 18144 5284
rect 17644 5244 17650 5256
rect 18138 5244 18144 5256
rect 18196 5284 18202 5296
rect 18196 5256 18276 5284
rect 18196 5244 18202 5256
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 9732 5188 10333 5216
rect 9732 5176 9738 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5216 11023 5219
rect 11146 5216 11152 5228
rect 11011 5188 11152 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11330 5216 11336 5228
rect 11291 5188 11336 5216
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12124 5188 12725 5216
rect 12124 5176 12130 5188
rect 12713 5185 12725 5188
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14366 5216 14372 5228
rect 14047 5188 14372 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 15102 5216 15108 5228
rect 15063 5188 15108 5216
rect 15102 5176 15108 5188
rect 15160 5216 15166 5228
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 15160 5188 16681 5216
rect 15160 5176 15166 5188
rect 16669 5185 16681 5188
rect 16715 5216 16727 5219
rect 17402 5216 17408 5228
rect 16715 5188 17408 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 18248 5225 18276 5256
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5216 18567 5219
rect 18598 5216 18604 5228
rect 18555 5188 18604 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19260 5216 19288 5312
rect 20254 5284 20260 5296
rect 20215 5256 20260 5284
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19260 5188 19809 5216
rect 19797 5185 19809 5188
rect 19843 5216 19855 5219
rect 20162 5216 20168 5228
rect 19843 5188 20168 5216
rect 19843 5185 19855 5188
rect 19797 5179 19855 5185
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 11112 5120 11253 5148
rect 11112 5108 11118 5120
rect 11241 5117 11253 5120
rect 11287 5148 11299 5151
rect 11514 5148 11520 5160
rect 11287 5120 11520 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 12986 5148 12992 5160
rect 12667 5120 12992 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 11146 5040 11152 5092
rect 11204 5080 11210 5092
rect 11698 5080 11704 5092
rect 11204 5052 11704 5080
rect 11204 5040 11210 5052
rect 11698 5040 11704 5052
rect 11756 5080 11762 5092
rect 12636 5080 12664 5111
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 16577 5151 16635 5157
rect 16577 5148 16589 5151
rect 16356 5120 16589 5148
rect 16356 5108 16362 5120
rect 16577 5117 16589 5120
rect 16623 5148 16635 5151
rect 17862 5148 17868 5160
rect 16623 5120 17868 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 17862 5108 17868 5120
rect 17920 5148 17926 5160
rect 18325 5151 18383 5157
rect 18325 5148 18337 5151
rect 17920 5120 18337 5148
rect 17920 5108 17926 5120
rect 18325 5117 18337 5120
rect 18371 5117 18383 5151
rect 18690 5148 18696 5160
rect 18651 5120 18696 5148
rect 18325 5111 18383 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 19150 5108 19156 5160
rect 19208 5148 19214 5160
rect 19705 5151 19763 5157
rect 19705 5148 19717 5151
rect 19208 5120 19717 5148
rect 19208 5108 19214 5120
rect 19705 5117 19717 5120
rect 19751 5148 19763 5151
rect 20438 5148 20444 5160
rect 19751 5120 20444 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 20438 5108 20444 5120
rect 20496 5148 20502 5160
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 20496 5120 21281 5148
rect 20496 5108 20502 5120
rect 21269 5117 21281 5120
rect 21315 5148 21327 5151
rect 21910 5148 21916 5160
rect 21315 5120 21916 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 11756 5052 12664 5080
rect 11756 5040 11762 5052
rect 8665 5015 8723 5021
rect 8665 4981 8677 5015
rect 8711 5012 8723 5015
rect 8754 5012 8760 5024
rect 8711 4984 8760 5012
rect 8711 4981 8723 4984
rect 8665 4975 8723 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9493 5015 9551 5021
rect 9493 4981 9505 5015
rect 9539 5012 9551 5015
rect 9674 5012 9680 5024
rect 9539 4984 9680 5012
rect 9539 4981 9551 4984
rect 9493 4975 9551 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 13630 5012 13636 5024
rect 13591 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 16390 4972 16396 5024
rect 16448 5012 16454 5024
rect 16853 5015 16911 5021
rect 16853 5012 16865 5015
rect 16448 4984 16865 5012
rect 16448 4972 16454 4984
rect 16853 4981 16865 4984
rect 16899 4981 16911 5015
rect 16853 4975 16911 4981
rect 1104 4922 28336 4944
rect 1104 4870 3282 4922
rect 3334 4870 3346 4922
rect 3398 4870 3410 4922
rect 3462 4870 3474 4922
rect 3526 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 6410 4922
rect 6462 4870 6474 4922
rect 6526 4870 9282 4922
rect 9334 4870 9346 4922
rect 9398 4870 9410 4922
rect 9462 4870 9474 4922
rect 9526 4870 12282 4922
rect 12334 4870 12346 4922
rect 12398 4870 12410 4922
rect 12462 4870 12474 4922
rect 12526 4870 15282 4922
rect 15334 4870 15346 4922
rect 15398 4870 15410 4922
rect 15462 4870 15474 4922
rect 15526 4870 18282 4922
rect 18334 4870 18346 4922
rect 18398 4870 18410 4922
rect 18462 4870 18474 4922
rect 18526 4870 21282 4922
rect 21334 4870 21346 4922
rect 21398 4870 21410 4922
rect 21462 4870 21474 4922
rect 21526 4870 24282 4922
rect 24334 4870 24346 4922
rect 24398 4870 24410 4922
rect 24462 4870 24474 4922
rect 24526 4870 27282 4922
rect 27334 4870 27346 4922
rect 27398 4870 27410 4922
rect 27462 4870 27474 4922
rect 27526 4870 28336 4922
rect 1104 4848 28336 4870
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 8110 4808 8116 4820
rect 7883 4780 8116 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 11054 4808 11060 4820
rect 8987 4780 11060 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 11054 4768 11060 4780
rect 11112 4808 11118 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 11112 4780 12633 4808
rect 11112 4768 11118 4780
rect 12621 4777 12633 4780
rect 12667 4808 12679 4811
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 12667 4780 13369 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 13357 4777 13369 4780
rect 13403 4808 13415 4811
rect 13630 4808 13636 4820
rect 13403 4780 13636 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14550 4808 14556 4820
rect 14511 4780 14556 4808
rect 14550 4768 14556 4780
rect 14608 4808 14614 4820
rect 18138 4808 18144 4820
rect 14608 4780 15424 4808
rect 18099 4780 18144 4808
rect 14608 4768 14614 4780
rect 15396 4752 15424 4780
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 19153 4811 19211 4817
rect 19153 4808 19165 4811
rect 18932 4780 19165 4808
rect 18932 4768 18938 4780
rect 19153 4777 19165 4780
rect 19199 4777 19211 4811
rect 19153 4771 19211 4777
rect 19610 4768 19616 4820
rect 19668 4808 19674 4820
rect 19889 4811 19947 4817
rect 19889 4808 19901 4811
rect 19668 4780 19901 4808
rect 19668 4768 19674 4780
rect 19889 4777 19901 4780
rect 19935 4777 19947 4811
rect 20162 4808 20168 4820
rect 20123 4780 20168 4808
rect 19889 4771 19947 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 8573 4743 8631 4749
rect 8573 4709 8585 4743
rect 8619 4740 8631 4743
rect 11330 4740 11336 4752
rect 8619 4712 11336 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 15378 4700 15384 4752
rect 15436 4700 15442 4752
rect 8202 4672 8208 4684
rect 8115 4644 8208 4672
rect 8202 4632 8208 4644
rect 8260 4672 8266 4684
rect 11422 4672 11428 4684
rect 8260 4644 11428 4672
rect 8260 4632 8266 4644
rect 11422 4632 11428 4644
rect 11480 4672 11486 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 11480 4644 11529 4672
rect 11480 4632 11486 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15160 4644 15485 4672
rect 15160 4632 15166 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 16114 4672 16120 4684
rect 16075 4644 16120 4672
rect 15473 4635 15531 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17862 4632 17868 4644
rect 17920 4672 17926 4684
rect 21085 4675 21143 4681
rect 21085 4672 21097 4675
rect 17920 4644 21097 4672
rect 17920 4632 17926 4644
rect 21085 4641 21097 4644
rect 21131 4672 21143 4675
rect 21453 4675 21511 4681
rect 21453 4672 21465 4675
rect 21131 4644 21465 4672
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 21453 4641 21465 4644
rect 21499 4641 21511 4675
rect 21453 4635 21511 4641
rect 10226 4604 10232 4616
rect 10139 4576 10232 4604
rect 10226 4564 10232 4576
rect 10284 4604 10290 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10284 4576 11069 4604
rect 10284 4564 10290 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 10410 4496 10416 4548
rect 10468 4536 10474 4548
rect 10505 4539 10563 4545
rect 10505 4536 10517 4539
rect 10468 4508 10517 4536
rect 10468 4496 10474 4508
rect 10505 4505 10517 4508
rect 10551 4505 10563 4539
rect 11348 4536 11376 4567
rect 11606 4564 11612 4616
rect 11664 4604 11670 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 11664 4576 13001 4604
rect 11664 4564 11670 4576
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 14182 4604 14188 4616
rect 13035 4576 14188 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 17218 4564 17224 4616
rect 17276 4564 17282 4616
rect 18138 4564 18144 4616
rect 18196 4604 18202 4616
rect 18598 4604 18604 4616
rect 18196 4576 18604 4604
rect 18196 4564 18202 4576
rect 18598 4564 18604 4576
rect 18656 4604 18662 4616
rect 18693 4607 18751 4613
rect 18693 4604 18705 4607
rect 18656 4576 18705 4604
rect 18656 4564 18662 4576
rect 18693 4573 18705 4576
rect 18739 4573 18751 4607
rect 18693 4567 18751 4573
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19668 4576 19717 4604
rect 19668 4564 19674 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 11882 4536 11888 4548
rect 11348 4508 11888 4536
rect 10505 4499 10563 4505
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 14921 4539 14979 4545
rect 13786 4508 14872 4536
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 8996 4440 9229 4468
rect 8996 4428 9002 4440
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 9217 4431 9275 4437
rect 11793 4471 11851 4477
rect 11793 4437 11805 4471
rect 11839 4468 11851 4471
rect 11974 4468 11980 4480
rect 11839 4440 11980 4468
rect 11839 4437 11851 4440
rect 11793 4431 11851 4437
rect 11974 4428 11980 4440
rect 12032 4468 12038 4480
rect 13786 4468 13814 4508
rect 12032 4440 13814 4468
rect 14093 4471 14151 4477
rect 12032 4428 12038 4440
rect 14093 4437 14105 4471
rect 14139 4468 14151 4471
rect 14366 4468 14372 4480
rect 14139 4440 14372 4468
rect 14139 4437 14151 4440
rect 14093 4431 14151 4437
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 14844 4468 14872 4508
rect 14921 4505 14933 4539
rect 14967 4536 14979 4539
rect 16390 4536 16396 4548
rect 14967 4508 16396 4536
rect 14967 4505 14979 4508
rect 14921 4499 14979 4505
rect 16390 4496 16396 4508
rect 16448 4496 16454 4548
rect 18782 4536 18788 4548
rect 17420 4508 18788 4536
rect 17420 4468 17448 4508
rect 18782 4496 18788 4508
rect 18840 4536 18846 4548
rect 18840 4508 18920 4536
rect 18840 4496 18846 4508
rect 18892 4477 18920 4508
rect 14844 4440 17448 4468
rect 18877 4471 18935 4477
rect 18877 4437 18889 4471
rect 18923 4437 18935 4471
rect 18877 4431 18935 4437
rect 1104 4378 28336 4400
rect 1104 4326 1782 4378
rect 1834 4326 1846 4378
rect 1898 4326 1910 4378
rect 1962 4326 1974 4378
rect 2026 4326 4782 4378
rect 4834 4326 4846 4378
rect 4898 4326 4910 4378
rect 4962 4326 4974 4378
rect 5026 4326 7782 4378
rect 7834 4326 7846 4378
rect 7898 4326 7910 4378
rect 7962 4326 7974 4378
rect 8026 4326 10782 4378
rect 10834 4326 10846 4378
rect 10898 4326 10910 4378
rect 10962 4326 10974 4378
rect 11026 4326 13782 4378
rect 13834 4326 13846 4378
rect 13898 4326 13910 4378
rect 13962 4326 13974 4378
rect 14026 4326 16782 4378
rect 16834 4326 16846 4378
rect 16898 4326 16910 4378
rect 16962 4326 16974 4378
rect 17026 4326 19782 4378
rect 19834 4326 19846 4378
rect 19898 4326 19910 4378
rect 19962 4326 19974 4378
rect 20026 4326 22782 4378
rect 22834 4326 22846 4378
rect 22898 4326 22910 4378
rect 22962 4326 22974 4378
rect 23026 4326 25782 4378
rect 25834 4326 25846 4378
rect 25898 4326 25910 4378
rect 25962 4326 25974 4378
rect 26026 4326 28336 4378
rect 1104 4304 28336 4326
rect 7837 4267 7895 4273
rect 7837 4233 7849 4267
rect 7883 4264 7895 4267
rect 8202 4264 8208 4276
rect 7883 4236 8208 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 14090 4264 14096 4276
rect 12676 4236 14096 4264
rect 12676 4224 12682 4236
rect 14090 4224 14096 4236
rect 14148 4264 14154 4276
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 14148 4236 15577 4264
rect 14148 4224 14154 4236
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 15565 4227 15623 4233
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19518 4264 19524 4276
rect 19383 4236 19524 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20438 4264 20444 4276
rect 20399 4236 20444 4264
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 9674 4196 9680 4208
rect 9171 4168 9680 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 9674 4156 9680 4168
rect 9732 4196 9738 4208
rect 9732 4168 10272 4196
rect 9732 4156 9738 4168
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11517 4199 11575 4205
rect 11517 4196 11529 4199
rect 11296 4168 11529 4196
rect 11296 4156 11302 4168
rect 11517 4165 11529 4168
rect 11563 4196 11575 4199
rect 11606 4196 11612 4208
rect 11563 4168 11612 4196
rect 11563 4165 11575 4168
rect 11517 4159 11575 4165
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 13538 4156 13544 4208
rect 13596 4196 13602 4208
rect 14458 4196 14464 4208
rect 13596 4168 14464 4196
rect 13596 4156 13602 4168
rect 14458 4156 14464 4168
rect 14516 4196 14522 4208
rect 16393 4199 16451 4205
rect 16393 4196 16405 4199
rect 14516 4168 16405 4196
rect 14516 4156 14522 4168
rect 16393 4165 16405 4168
rect 16439 4196 16451 4199
rect 16666 4196 16672 4208
rect 16439 4168 16672 4196
rect 16439 4165 16451 4168
rect 16393 4159 16451 4165
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 8110 4128 8116 4140
rect 8071 4100 8116 4128
rect 8110 4088 8116 4100
rect 8168 4088 8174 4140
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8754 4128 8760 4140
rect 8343 4100 8760 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 8312 4060 8340 4091
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 15378 4128 15384 4140
rect 15339 4100 15384 4128
rect 14001 4091 14059 4097
rect 8662 4060 8668 4072
rect 7515 4032 8340 4060
rect 8623 4032 8668 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 9122 4060 9128 4072
rect 8904 4032 9128 4060
rect 8904 4020 8910 4032
rect 9122 4020 9128 4032
rect 9180 4060 9186 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9180 4032 9505 4060
rect 9180 4020 9186 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9766 4060 9772 4072
rect 9727 4032 9772 4060
rect 9493 4023 9551 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 11238 4060 11244 4072
rect 10192 4032 11244 4060
rect 10192 4020 10198 4032
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 14016 3992 14044 4091
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 18138 4128 18144 4140
rect 17083 4100 18144 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 18690 4128 18696 4140
rect 18651 4100 18696 4128
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 19610 4128 19616 4140
rect 19571 4100 19616 4128
rect 19610 4088 19616 4100
rect 19668 4128 19674 4140
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19668 4100 20085 4128
rect 19668 4088 19674 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 14148 4032 18245 4060
rect 14148 4020 14154 4032
rect 18233 4029 18245 4032
rect 18279 4029 18291 4063
rect 18233 4023 18291 4029
rect 15105 3995 15163 4001
rect 14016 3964 14504 3992
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 11296 3896 12909 3924
rect 11296 3884 11302 3896
rect 12897 3893 12909 3896
rect 12943 3924 12955 3927
rect 13170 3924 13176 3936
rect 12943 3896 13176 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13170 3884 13176 3896
rect 13228 3924 13234 3936
rect 13630 3924 13636 3936
rect 13228 3896 13636 3924
rect 13228 3884 13234 3896
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 14476 3933 14504 3964
rect 15105 3961 15117 3995
rect 15151 3992 15163 3995
rect 17218 3992 17224 4004
rect 15151 3964 17224 3992
rect 15151 3961 15163 3964
rect 15105 3955 15163 3961
rect 17218 3952 17224 3964
rect 17276 3992 17282 4004
rect 19797 3995 19855 4001
rect 19797 3992 19809 3995
rect 17276 3964 19809 3992
rect 17276 3952 17282 3964
rect 19797 3961 19809 3964
rect 19843 3961 19855 3995
rect 19797 3955 19855 3961
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 15010 3924 15016 3936
rect 14507 3896 15016 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 15010 3884 15016 3896
rect 15068 3884 15074 3936
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 15933 3927 15991 3933
rect 15933 3924 15945 3927
rect 15896 3896 15945 3924
rect 15896 3884 15902 3896
rect 15933 3893 15945 3896
rect 15979 3924 15991 3927
rect 16206 3924 16212 3936
rect 15979 3896 16212 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 1104 3834 28336 3856
rect 1104 3782 3282 3834
rect 3334 3782 3346 3834
rect 3398 3782 3410 3834
rect 3462 3782 3474 3834
rect 3526 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 6410 3834
rect 6462 3782 6474 3834
rect 6526 3782 9282 3834
rect 9334 3782 9346 3834
rect 9398 3782 9410 3834
rect 9462 3782 9474 3834
rect 9526 3782 12282 3834
rect 12334 3782 12346 3834
rect 12398 3782 12410 3834
rect 12462 3782 12474 3834
rect 12526 3782 15282 3834
rect 15334 3782 15346 3834
rect 15398 3782 15410 3834
rect 15462 3782 15474 3834
rect 15526 3782 18282 3834
rect 18334 3782 18346 3834
rect 18398 3782 18410 3834
rect 18462 3782 18474 3834
rect 18526 3782 21282 3834
rect 21334 3782 21346 3834
rect 21398 3782 21410 3834
rect 21462 3782 21474 3834
rect 21526 3782 24282 3834
rect 24334 3782 24346 3834
rect 24398 3782 24410 3834
rect 24462 3782 24474 3834
rect 24526 3782 27282 3834
rect 27334 3782 27346 3834
rect 27398 3782 27410 3834
rect 27462 3782 27474 3834
rect 27526 3782 28336 3834
rect 1104 3760 28336 3782
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 8754 3720 8760 3732
rect 8619 3692 8760 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 10226 3720 10232 3732
rect 9692 3692 10232 3720
rect 8110 3612 8116 3664
rect 8168 3652 8174 3664
rect 8205 3655 8263 3661
rect 8205 3652 8217 3655
rect 8168 3624 8217 3652
rect 8168 3612 8174 3624
rect 8205 3621 8217 3624
rect 8251 3652 8263 3655
rect 9692 3652 9720 3692
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12713 3723 12771 3729
rect 12713 3720 12725 3723
rect 11940 3692 12725 3720
rect 11940 3680 11946 3692
rect 12713 3689 12725 3692
rect 12759 3689 12771 3723
rect 12713 3683 12771 3689
rect 8251 3624 9720 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 12728 3516 12756 3683
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 14461 3723 14519 3729
rect 14461 3720 14473 3723
rect 13688 3692 14473 3720
rect 13688 3680 13694 3692
rect 14461 3689 14473 3692
rect 14507 3689 14519 3723
rect 14461 3683 14519 3689
rect 15933 3723 15991 3729
rect 15933 3689 15945 3723
rect 15979 3720 15991 3723
rect 16114 3720 16120 3732
rect 15979 3692 16120 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 18785 3723 18843 3729
rect 18785 3720 18797 3723
rect 18748 3692 18797 3720
rect 18748 3680 18754 3692
rect 18785 3689 18797 3692
rect 18831 3689 18843 3723
rect 18785 3683 18843 3689
rect 15562 3652 15568 3664
rect 15523 3624 15568 3652
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 14090 3584 14096 3596
rect 14051 3556 14096 3584
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3584 16819 3587
rect 17218 3584 17224 3596
rect 16807 3556 17224 3584
rect 16807 3553 16819 3556
rect 16761 3547 16819 3553
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3584 18202 3596
rect 19058 3584 19064 3596
rect 18196 3556 19064 3584
rect 18196 3544 18202 3556
rect 19058 3544 19064 3556
rect 19116 3584 19122 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 19116 3556 19165 3584
rect 19116 3544 19122 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19153 3547 19211 3553
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12728 3488 13093 3516
rect 10137 3479 10195 3485
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13081 3479 13139 3485
rect 8941 3451 8999 3457
rect 8941 3417 8953 3451
rect 8987 3448 8999 3451
rect 9766 3448 9772 3460
rect 8987 3420 9772 3448
rect 8987 3417 8999 3420
rect 8941 3411 8999 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 9180 3352 9229 3380
rect 9180 3340 9186 3352
rect 9217 3349 9229 3352
rect 9263 3380 9275 3383
rect 10152 3380 10180 3479
rect 10410 3448 10416 3460
rect 10371 3420 10416 3448
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 10502 3408 10508 3460
rect 10560 3448 10566 3460
rect 12158 3448 12164 3460
rect 10560 3420 10916 3448
rect 12119 3420 12164 3448
rect 10560 3408 10566 3420
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 13096 3448 13124 3479
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 16206 3476 16212 3528
rect 16264 3516 16270 3528
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 16264 3488 16405 3516
rect 16264 3476 16270 3488
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 19610 3516 19616 3528
rect 18656 3488 19616 3516
rect 18656 3476 18662 3488
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 16298 3448 16304 3460
rect 13096 3420 16304 3448
rect 16298 3408 16304 3420
rect 16356 3408 16362 3460
rect 17770 3408 17776 3460
rect 17828 3408 17834 3460
rect 13170 3380 13176 3392
rect 9263 3352 10180 3380
rect 13131 3352 13176 3380
rect 9263 3349 9275 3352
rect 9217 3343 9275 3349
rect 13170 3340 13176 3352
rect 13228 3340 13234 3392
rect 14921 3383 14979 3389
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 15010 3380 15016 3392
rect 14967 3352 15016 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 1104 3290 28336 3312
rect 1104 3238 1782 3290
rect 1834 3238 1846 3290
rect 1898 3238 1910 3290
rect 1962 3238 1974 3290
rect 2026 3238 4782 3290
rect 4834 3238 4846 3290
rect 4898 3238 4910 3290
rect 4962 3238 4974 3290
rect 5026 3238 7782 3290
rect 7834 3238 7846 3290
rect 7898 3238 7910 3290
rect 7962 3238 7974 3290
rect 8026 3238 10782 3290
rect 10834 3238 10846 3290
rect 10898 3238 10910 3290
rect 10962 3238 10974 3290
rect 11026 3238 13782 3290
rect 13834 3238 13846 3290
rect 13898 3238 13910 3290
rect 13962 3238 13974 3290
rect 14026 3238 16782 3290
rect 16834 3238 16846 3290
rect 16898 3238 16910 3290
rect 16962 3238 16974 3290
rect 17026 3238 19782 3290
rect 19834 3238 19846 3290
rect 19898 3238 19910 3290
rect 19962 3238 19974 3290
rect 20026 3238 22782 3290
rect 22834 3238 22846 3290
rect 22898 3238 22910 3290
rect 22962 3238 22974 3290
rect 23026 3238 25782 3290
rect 25834 3238 25846 3290
rect 25898 3238 25910 3290
rect 25962 3238 25974 3290
rect 26026 3238 28336 3290
rect 1104 3216 28336 3238
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 8849 3179 8907 3185
rect 8849 3176 8861 3179
rect 8812 3148 8861 3176
rect 8812 3136 8818 3148
rect 8849 3145 8861 3148
rect 8895 3145 8907 3179
rect 8849 3139 8907 3145
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 12066 3176 12072 3188
rect 11011 3148 12072 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12805 3179 12863 3185
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 12851 3148 14504 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 14476 3120 14504 3148
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 17405 3139 17463 3145
rect 19058 3136 19064 3148
rect 19116 3176 19122 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 19116 3148 19441 3176
rect 19116 3136 19122 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 19429 3139 19487 3145
rect 9766 3108 9772 3120
rect 9727 3080 9772 3108
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 10226 3068 10232 3120
rect 10284 3108 10290 3120
rect 10284 3080 10640 3108
rect 10284 3068 10290 3080
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 8720 3012 9689 3040
rect 8720 3000 8726 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10612 3049 10640 3080
rect 13170 3068 13176 3120
rect 13228 3108 13234 3120
rect 14001 3111 14059 3117
rect 14001 3108 14013 3111
rect 13228 3080 14013 3108
rect 13228 3068 13234 3080
rect 14001 3077 14013 3080
rect 14047 3077 14059 3111
rect 14001 3071 14059 3077
rect 14458 3068 14464 3120
rect 14516 3068 14522 3120
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10192 3012 10517 3040
rect 10192 3000 10198 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3040 10655 3043
rect 11330 3040 11336 3052
rect 10643 3012 11336 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 12618 3040 12624 3052
rect 12575 3012 12624 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18196 3012 18245 3040
rect 18196 3000 18202 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11425 2975 11483 2981
rect 11425 2972 11437 2975
rect 11020 2944 11437 2972
rect 11020 2932 11026 2944
rect 11425 2941 11437 2944
rect 11471 2972 11483 2975
rect 13722 2972 13728 2984
rect 11471 2944 13216 2972
rect 13683 2944 13728 2972
rect 11471 2941 11483 2944
rect 11425 2935 11483 2941
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 13188 2913 13216 2944
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14090 2972 14096 2984
rect 13832 2944 14096 2972
rect 11977 2907 12035 2913
rect 11977 2904 11989 2907
rect 10836 2876 11989 2904
rect 10836 2864 10842 2876
rect 11977 2873 11989 2876
rect 12023 2904 12035 2907
rect 12529 2907 12587 2913
rect 12529 2904 12541 2907
rect 12023 2876 12541 2904
rect 12023 2873 12035 2876
rect 11977 2867 12035 2873
rect 12529 2873 12541 2876
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 13173 2907 13231 2913
rect 13173 2873 13185 2907
rect 13219 2904 13231 2907
rect 13832 2904 13860 2944
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 15068 2944 15761 2972
rect 15068 2932 15074 2944
rect 15749 2941 15761 2944
rect 15795 2972 15807 2975
rect 16577 2975 16635 2981
rect 16577 2972 16589 2975
rect 15795 2944 16589 2972
rect 15795 2941 15807 2944
rect 15749 2935 15807 2941
rect 16577 2941 16589 2944
rect 16623 2972 16635 2975
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 16623 2944 18705 2972
rect 16623 2941 16635 2944
rect 16577 2935 16635 2941
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 18693 2935 18751 2941
rect 13219 2876 13860 2904
rect 13219 2873 13231 2876
rect 13173 2867 13231 2873
rect 15562 2864 15568 2916
rect 15620 2904 15626 2916
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 15620 2876 18429 2904
rect 15620 2864 15626 2876
rect 18417 2873 18429 2876
rect 18463 2904 18475 2907
rect 18598 2904 18604 2916
rect 18463 2876 18604 2904
rect 18463 2873 18475 2876
rect 18417 2867 18475 2873
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 10502 2836 10508 2848
rect 9355 2808 10508 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 16206 2836 16212 2848
rect 13780 2808 16212 2836
rect 13780 2796 13786 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 16356 2808 16865 2836
rect 16356 2796 16362 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 1104 2746 28336 2768
rect 1104 2694 3282 2746
rect 3334 2694 3346 2746
rect 3398 2694 3410 2746
rect 3462 2694 3474 2746
rect 3526 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 6410 2746
rect 6462 2694 6474 2746
rect 6526 2694 9282 2746
rect 9334 2694 9346 2746
rect 9398 2694 9410 2746
rect 9462 2694 9474 2746
rect 9526 2694 12282 2746
rect 12334 2694 12346 2746
rect 12398 2694 12410 2746
rect 12462 2694 12474 2746
rect 12526 2694 15282 2746
rect 15334 2694 15346 2746
rect 15398 2694 15410 2746
rect 15462 2694 15474 2746
rect 15526 2694 18282 2746
rect 18334 2694 18346 2746
rect 18398 2694 18410 2746
rect 18462 2694 18474 2746
rect 18526 2694 21282 2746
rect 21334 2694 21346 2746
rect 21398 2694 21410 2746
rect 21462 2694 21474 2746
rect 21526 2694 24282 2746
rect 24334 2694 24346 2746
rect 24398 2694 24410 2746
rect 24462 2694 24474 2746
rect 24526 2694 27282 2746
rect 27334 2694 27346 2746
rect 27398 2694 27410 2746
rect 27462 2694 27474 2746
rect 27526 2694 28336 2746
rect 1104 2672 28336 2694
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8720 2604 8953 2632
rect 8720 2592 8726 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10502 2632 10508 2644
rect 10183 2604 10508 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 13170 2632 13176 2644
rect 13131 2604 13176 2632
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14516 2604 14841 2632
rect 14516 2592 14522 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 16025 2635 16083 2641
rect 16025 2601 16037 2635
rect 16071 2632 16083 2635
rect 17770 2632 17776 2644
rect 16071 2604 17776 2632
rect 16071 2601 16083 2604
rect 16025 2595 16083 2601
rect 17770 2592 17776 2604
rect 17828 2632 17834 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 17828 2604 18705 2632
rect 17828 2592 17834 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 10410 2564 10416 2576
rect 10371 2536 10416 2564
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 12253 2567 12311 2573
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 13538 2564 13544 2576
rect 12299 2536 13544 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 13538 2524 13544 2536
rect 13596 2564 13602 2576
rect 13955 2567 14013 2573
rect 13955 2564 13967 2567
rect 13596 2536 13967 2564
rect 13596 2524 13602 2536
rect 13955 2533 13967 2536
rect 14001 2533 14013 2567
rect 13955 2527 14013 2533
rect 14093 2567 14151 2573
rect 14093 2533 14105 2567
rect 14139 2564 14151 2567
rect 19705 2567 19763 2573
rect 19705 2564 19717 2567
rect 14139 2536 19717 2564
rect 14139 2533 14151 2536
rect 14093 2527 14151 2533
rect 19705 2533 19717 2536
rect 19751 2533 19763 2567
rect 19705 2527 19763 2533
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2496 7987 2499
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 7975 2468 11069 2496
rect 7975 2465 7987 2468
rect 7929 2459 7987 2465
rect 11057 2465 11069 2468
rect 11103 2496 11115 2499
rect 11146 2496 11152 2508
rect 11103 2468 11152 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 11146 2456 11152 2468
rect 11204 2456 11210 2508
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11388 2468 11437 2496
rect 11388 2456 11394 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 14108 2496 14136 2527
rect 12216 2468 14136 2496
rect 14185 2499 14243 2505
rect 12216 2456 12222 2468
rect 14185 2465 14197 2499
rect 14231 2496 14243 2499
rect 15010 2496 15016 2508
rect 14231 2468 15016 2496
rect 14231 2465 14243 2468
rect 14185 2459 14243 2465
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 17773 2499 17831 2505
rect 17773 2496 17785 2499
rect 16724 2468 17785 2496
rect 16724 2456 16730 2468
rect 17773 2465 17785 2468
rect 17819 2496 17831 2499
rect 18690 2496 18696 2508
rect 17819 2468 18696 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 8938 2428 8944 2440
rect 8711 2400 8944 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 8938 2388 8944 2400
rect 8996 2428 9002 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 8996 2400 9965 2428
rect 8996 2388 9002 2400
rect 9953 2397 9965 2400
rect 9999 2428 10011 2431
rect 10778 2428 10784 2440
rect 9999 2400 10784 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11238 2428 11244 2440
rect 11199 2400 11244 2428
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 9401 2363 9459 2369
rect 9401 2329 9413 2363
rect 9447 2360 9459 2363
rect 11348 2360 11376 2456
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 12124 2400 13461 2428
rect 12124 2388 12130 2400
rect 13449 2397 13461 2400
rect 13495 2428 13507 2431
rect 13722 2428 13728 2440
rect 13495 2400 13728 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 16393 2431 16451 2437
rect 16393 2397 16405 2431
rect 16439 2428 16451 2431
rect 17313 2431 17371 2437
rect 17313 2428 17325 2431
rect 16439 2400 17325 2428
rect 16439 2397 16451 2400
rect 16393 2391 16451 2397
rect 17313 2397 17325 2400
rect 17359 2428 17371 2431
rect 18230 2428 18236 2440
rect 17359 2400 18236 2428
rect 17359 2397 17371 2400
rect 17313 2391 17371 2397
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 18509 2431 18567 2437
rect 18509 2397 18521 2431
rect 18555 2428 18567 2431
rect 18598 2428 18604 2440
rect 18555 2400 18604 2428
rect 18555 2397 18567 2400
rect 18509 2391 18567 2397
rect 18598 2388 18604 2400
rect 18656 2428 18662 2440
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 18656 2400 19349 2428
rect 18656 2388 18662 2400
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 19337 2391 19395 2397
rect 9447 2332 11376 2360
rect 13817 2363 13875 2369
rect 9447 2329 9459 2332
rect 9401 2323 9459 2329
rect 13817 2329 13829 2363
rect 13863 2329 13875 2363
rect 13817 2323 13875 2329
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 11238 2292 11244 2304
rect 8343 2264 11244 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 13832 2292 13860 2323
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 16669 2363 16727 2369
rect 16669 2360 16681 2363
rect 14424 2332 16681 2360
rect 14424 2320 14430 2332
rect 16669 2329 16681 2332
rect 16715 2360 16727 2363
rect 18138 2360 18144 2372
rect 16715 2332 18144 2360
rect 16715 2329 16727 2332
rect 16669 2323 16727 2329
rect 18138 2320 18144 2332
rect 18196 2360 18202 2372
rect 18969 2363 19027 2369
rect 18969 2360 18981 2363
rect 18196 2332 18981 2360
rect 18196 2320 18202 2332
rect 18969 2329 18981 2332
rect 19015 2329 19027 2363
rect 18969 2323 19027 2329
rect 14182 2292 14188 2304
rect 13832 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2292 14246 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 14240 2264 20085 2292
rect 14240 2252 14246 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 1104 2202 28336 2224
rect 1104 2150 1782 2202
rect 1834 2150 1846 2202
rect 1898 2150 1910 2202
rect 1962 2150 1974 2202
rect 2026 2150 4782 2202
rect 4834 2150 4846 2202
rect 4898 2150 4910 2202
rect 4962 2150 4974 2202
rect 5026 2150 7782 2202
rect 7834 2150 7846 2202
rect 7898 2150 7910 2202
rect 7962 2150 7974 2202
rect 8026 2150 10782 2202
rect 10834 2150 10846 2202
rect 10898 2150 10910 2202
rect 10962 2150 10974 2202
rect 11026 2150 13782 2202
rect 13834 2150 13846 2202
rect 13898 2150 13910 2202
rect 13962 2150 13974 2202
rect 14026 2150 16782 2202
rect 16834 2150 16846 2202
rect 16898 2150 16910 2202
rect 16962 2150 16974 2202
rect 17026 2150 19782 2202
rect 19834 2150 19846 2202
rect 19898 2150 19910 2202
rect 19962 2150 19974 2202
rect 20026 2150 22782 2202
rect 22834 2150 22846 2202
rect 22898 2150 22910 2202
rect 22962 2150 22974 2202
rect 23026 2150 25782 2202
rect 25834 2150 25846 2202
rect 25898 2150 25910 2202
rect 25962 2150 25974 2202
rect 26026 2150 28336 2202
rect 1104 2128 28336 2150
rect 290 1300 296 1352
rect 348 1340 354 1352
rect 10318 1340 10324 1352
rect 348 1312 10324 1340
rect 348 1300 354 1312
rect 10318 1300 10324 1312
rect 10376 1300 10382 1352
<< via1 >>
rect 1782 29350 1834 29402
rect 1846 29350 1898 29402
rect 1910 29350 1962 29402
rect 1974 29350 2026 29402
rect 4782 29350 4834 29402
rect 4846 29350 4898 29402
rect 4910 29350 4962 29402
rect 4974 29350 5026 29402
rect 7782 29350 7834 29402
rect 7846 29350 7898 29402
rect 7910 29350 7962 29402
rect 7974 29350 8026 29402
rect 10782 29350 10834 29402
rect 10846 29350 10898 29402
rect 10910 29350 10962 29402
rect 10974 29350 11026 29402
rect 13782 29350 13834 29402
rect 13846 29350 13898 29402
rect 13910 29350 13962 29402
rect 13974 29350 14026 29402
rect 16782 29350 16834 29402
rect 16846 29350 16898 29402
rect 16910 29350 16962 29402
rect 16974 29350 17026 29402
rect 19782 29350 19834 29402
rect 19846 29350 19898 29402
rect 19910 29350 19962 29402
rect 19974 29350 20026 29402
rect 22782 29350 22834 29402
rect 22846 29350 22898 29402
rect 22910 29350 22962 29402
rect 22974 29350 23026 29402
rect 25782 29350 25834 29402
rect 25846 29350 25898 29402
rect 25910 29350 25962 29402
rect 25974 29350 26026 29402
rect 3282 28806 3334 28858
rect 3346 28806 3398 28858
rect 3410 28806 3462 28858
rect 3474 28806 3526 28858
rect 6282 28806 6334 28858
rect 6346 28806 6398 28858
rect 6410 28806 6462 28858
rect 6474 28806 6526 28858
rect 9282 28806 9334 28858
rect 9346 28806 9398 28858
rect 9410 28806 9462 28858
rect 9474 28806 9526 28858
rect 12282 28806 12334 28858
rect 12346 28806 12398 28858
rect 12410 28806 12462 28858
rect 12474 28806 12526 28858
rect 15282 28806 15334 28858
rect 15346 28806 15398 28858
rect 15410 28806 15462 28858
rect 15474 28806 15526 28858
rect 18282 28806 18334 28858
rect 18346 28806 18398 28858
rect 18410 28806 18462 28858
rect 18474 28806 18526 28858
rect 21282 28806 21334 28858
rect 21346 28806 21398 28858
rect 21410 28806 21462 28858
rect 21474 28806 21526 28858
rect 24282 28806 24334 28858
rect 24346 28806 24398 28858
rect 24410 28806 24462 28858
rect 24474 28806 24526 28858
rect 27282 28806 27334 28858
rect 27346 28806 27398 28858
rect 27410 28806 27462 28858
rect 27474 28806 27526 28858
rect 1782 28262 1834 28314
rect 1846 28262 1898 28314
rect 1910 28262 1962 28314
rect 1974 28262 2026 28314
rect 4782 28262 4834 28314
rect 4846 28262 4898 28314
rect 4910 28262 4962 28314
rect 4974 28262 5026 28314
rect 7782 28262 7834 28314
rect 7846 28262 7898 28314
rect 7910 28262 7962 28314
rect 7974 28262 8026 28314
rect 10782 28262 10834 28314
rect 10846 28262 10898 28314
rect 10910 28262 10962 28314
rect 10974 28262 11026 28314
rect 13782 28262 13834 28314
rect 13846 28262 13898 28314
rect 13910 28262 13962 28314
rect 13974 28262 14026 28314
rect 16782 28262 16834 28314
rect 16846 28262 16898 28314
rect 16910 28262 16962 28314
rect 16974 28262 17026 28314
rect 19782 28262 19834 28314
rect 19846 28262 19898 28314
rect 19910 28262 19962 28314
rect 19974 28262 20026 28314
rect 22782 28262 22834 28314
rect 22846 28262 22898 28314
rect 22910 28262 22962 28314
rect 22974 28262 23026 28314
rect 25782 28262 25834 28314
rect 25846 28262 25898 28314
rect 25910 28262 25962 28314
rect 25974 28262 26026 28314
rect 3282 27718 3334 27770
rect 3346 27718 3398 27770
rect 3410 27718 3462 27770
rect 3474 27718 3526 27770
rect 6282 27718 6334 27770
rect 6346 27718 6398 27770
rect 6410 27718 6462 27770
rect 6474 27718 6526 27770
rect 9282 27718 9334 27770
rect 9346 27718 9398 27770
rect 9410 27718 9462 27770
rect 9474 27718 9526 27770
rect 12282 27718 12334 27770
rect 12346 27718 12398 27770
rect 12410 27718 12462 27770
rect 12474 27718 12526 27770
rect 15282 27718 15334 27770
rect 15346 27718 15398 27770
rect 15410 27718 15462 27770
rect 15474 27718 15526 27770
rect 18282 27718 18334 27770
rect 18346 27718 18398 27770
rect 18410 27718 18462 27770
rect 18474 27718 18526 27770
rect 21282 27718 21334 27770
rect 21346 27718 21398 27770
rect 21410 27718 21462 27770
rect 21474 27718 21526 27770
rect 24282 27718 24334 27770
rect 24346 27718 24398 27770
rect 24410 27718 24462 27770
rect 24474 27718 24526 27770
rect 27282 27718 27334 27770
rect 27346 27718 27398 27770
rect 27410 27718 27462 27770
rect 27474 27718 27526 27770
rect 23204 27412 23256 27464
rect 24584 27412 24636 27464
rect 23112 27387 23164 27396
rect 23112 27353 23121 27387
rect 23121 27353 23155 27387
rect 23155 27353 23164 27387
rect 23112 27344 23164 27353
rect 1782 27174 1834 27226
rect 1846 27174 1898 27226
rect 1910 27174 1962 27226
rect 1974 27174 2026 27226
rect 4782 27174 4834 27226
rect 4846 27174 4898 27226
rect 4910 27174 4962 27226
rect 4974 27174 5026 27226
rect 7782 27174 7834 27226
rect 7846 27174 7898 27226
rect 7910 27174 7962 27226
rect 7974 27174 8026 27226
rect 10782 27174 10834 27226
rect 10846 27174 10898 27226
rect 10910 27174 10962 27226
rect 10974 27174 11026 27226
rect 13782 27174 13834 27226
rect 13846 27174 13898 27226
rect 13910 27174 13962 27226
rect 13974 27174 14026 27226
rect 16782 27174 16834 27226
rect 16846 27174 16898 27226
rect 16910 27174 16962 27226
rect 16974 27174 17026 27226
rect 19782 27174 19834 27226
rect 19846 27174 19898 27226
rect 19910 27174 19962 27226
rect 19974 27174 20026 27226
rect 22782 27174 22834 27226
rect 22846 27174 22898 27226
rect 22910 27174 22962 27226
rect 22974 27174 23026 27226
rect 25782 27174 25834 27226
rect 25846 27174 25898 27226
rect 25910 27174 25962 27226
rect 25974 27174 26026 27226
rect 23204 27115 23256 27124
rect 23204 27081 23213 27115
rect 23213 27081 23247 27115
rect 23247 27081 23256 27115
rect 23204 27072 23256 27081
rect 3282 26630 3334 26682
rect 3346 26630 3398 26682
rect 3410 26630 3462 26682
rect 3474 26630 3526 26682
rect 6282 26630 6334 26682
rect 6346 26630 6398 26682
rect 6410 26630 6462 26682
rect 6474 26630 6526 26682
rect 9282 26630 9334 26682
rect 9346 26630 9398 26682
rect 9410 26630 9462 26682
rect 9474 26630 9526 26682
rect 12282 26630 12334 26682
rect 12346 26630 12398 26682
rect 12410 26630 12462 26682
rect 12474 26630 12526 26682
rect 15282 26630 15334 26682
rect 15346 26630 15398 26682
rect 15410 26630 15462 26682
rect 15474 26630 15526 26682
rect 18282 26630 18334 26682
rect 18346 26630 18398 26682
rect 18410 26630 18462 26682
rect 18474 26630 18526 26682
rect 21282 26630 21334 26682
rect 21346 26630 21398 26682
rect 21410 26630 21462 26682
rect 21474 26630 21526 26682
rect 24282 26630 24334 26682
rect 24346 26630 24398 26682
rect 24410 26630 24462 26682
rect 24474 26630 24526 26682
rect 27282 26630 27334 26682
rect 27346 26630 27398 26682
rect 27410 26630 27462 26682
rect 27474 26630 27526 26682
rect 1782 26086 1834 26138
rect 1846 26086 1898 26138
rect 1910 26086 1962 26138
rect 1974 26086 2026 26138
rect 4782 26086 4834 26138
rect 4846 26086 4898 26138
rect 4910 26086 4962 26138
rect 4974 26086 5026 26138
rect 7782 26086 7834 26138
rect 7846 26086 7898 26138
rect 7910 26086 7962 26138
rect 7974 26086 8026 26138
rect 10782 26086 10834 26138
rect 10846 26086 10898 26138
rect 10910 26086 10962 26138
rect 10974 26086 11026 26138
rect 13782 26086 13834 26138
rect 13846 26086 13898 26138
rect 13910 26086 13962 26138
rect 13974 26086 14026 26138
rect 16782 26086 16834 26138
rect 16846 26086 16898 26138
rect 16910 26086 16962 26138
rect 16974 26086 17026 26138
rect 19782 26086 19834 26138
rect 19846 26086 19898 26138
rect 19910 26086 19962 26138
rect 19974 26086 20026 26138
rect 22782 26086 22834 26138
rect 22846 26086 22898 26138
rect 22910 26086 22962 26138
rect 22974 26086 23026 26138
rect 25782 26086 25834 26138
rect 25846 26086 25898 26138
rect 25910 26086 25962 26138
rect 25974 26086 26026 26138
rect 3282 25542 3334 25594
rect 3346 25542 3398 25594
rect 3410 25542 3462 25594
rect 3474 25542 3526 25594
rect 6282 25542 6334 25594
rect 6346 25542 6398 25594
rect 6410 25542 6462 25594
rect 6474 25542 6526 25594
rect 9282 25542 9334 25594
rect 9346 25542 9398 25594
rect 9410 25542 9462 25594
rect 9474 25542 9526 25594
rect 12282 25542 12334 25594
rect 12346 25542 12398 25594
rect 12410 25542 12462 25594
rect 12474 25542 12526 25594
rect 15282 25542 15334 25594
rect 15346 25542 15398 25594
rect 15410 25542 15462 25594
rect 15474 25542 15526 25594
rect 18282 25542 18334 25594
rect 18346 25542 18398 25594
rect 18410 25542 18462 25594
rect 18474 25542 18526 25594
rect 21282 25542 21334 25594
rect 21346 25542 21398 25594
rect 21410 25542 21462 25594
rect 21474 25542 21526 25594
rect 24282 25542 24334 25594
rect 24346 25542 24398 25594
rect 24410 25542 24462 25594
rect 24474 25542 24526 25594
rect 27282 25542 27334 25594
rect 27346 25542 27398 25594
rect 27410 25542 27462 25594
rect 27474 25542 27526 25594
rect 1782 24998 1834 25050
rect 1846 24998 1898 25050
rect 1910 24998 1962 25050
rect 1974 24998 2026 25050
rect 4782 24998 4834 25050
rect 4846 24998 4898 25050
rect 4910 24998 4962 25050
rect 4974 24998 5026 25050
rect 7782 24998 7834 25050
rect 7846 24998 7898 25050
rect 7910 24998 7962 25050
rect 7974 24998 8026 25050
rect 10782 24998 10834 25050
rect 10846 24998 10898 25050
rect 10910 24998 10962 25050
rect 10974 24998 11026 25050
rect 13782 24998 13834 25050
rect 13846 24998 13898 25050
rect 13910 24998 13962 25050
rect 13974 24998 14026 25050
rect 16782 24998 16834 25050
rect 16846 24998 16898 25050
rect 16910 24998 16962 25050
rect 16974 24998 17026 25050
rect 19782 24998 19834 25050
rect 19846 24998 19898 25050
rect 19910 24998 19962 25050
rect 19974 24998 20026 25050
rect 22782 24998 22834 25050
rect 22846 24998 22898 25050
rect 22910 24998 22962 25050
rect 22974 24998 23026 25050
rect 25782 24998 25834 25050
rect 25846 24998 25898 25050
rect 25910 24998 25962 25050
rect 25974 24998 26026 25050
rect 3282 24454 3334 24506
rect 3346 24454 3398 24506
rect 3410 24454 3462 24506
rect 3474 24454 3526 24506
rect 6282 24454 6334 24506
rect 6346 24454 6398 24506
rect 6410 24454 6462 24506
rect 6474 24454 6526 24506
rect 9282 24454 9334 24506
rect 9346 24454 9398 24506
rect 9410 24454 9462 24506
rect 9474 24454 9526 24506
rect 12282 24454 12334 24506
rect 12346 24454 12398 24506
rect 12410 24454 12462 24506
rect 12474 24454 12526 24506
rect 15282 24454 15334 24506
rect 15346 24454 15398 24506
rect 15410 24454 15462 24506
rect 15474 24454 15526 24506
rect 18282 24454 18334 24506
rect 18346 24454 18398 24506
rect 18410 24454 18462 24506
rect 18474 24454 18526 24506
rect 21282 24454 21334 24506
rect 21346 24454 21398 24506
rect 21410 24454 21462 24506
rect 21474 24454 21526 24506
rect 24282 24454 24334 24506
rect 24346 24454 24398 24506
rect 24410 24454 24462 24506
rect 24474 24454 24526 24506
rect 27282 24454 27334 24506
rect 27346 24454 27398 24506
rect 27410 24454 27462 24506
rect 27474 24454 27526 24506
rect 1782 23910 1834 23962
rect 1846 23910 1898 23962
rect 1910 23910 1962 23962
rect 1974 23910 2026 23962
rect 4782 23910 4834 23962
rect 4846 23910 4898 23962
rect 4910 23910 4962 23962
rect 4974 23910 5026 23962
rect 7782 23910 7834 23962
rect 7846 23910 7898 23962
rect 7910 23910 7962 23962
rect 7974 23910 8026 23962
rect 10782 23910 10834 23962
rect 10846 23910 10898 23962
rect 10910 23910 10962 23962
rect 10974 23910 11026 23962
rect 13782 23910 13834 23962
rect 13846 23910 13898 23962
rect 13910 23910 13962 23962
rect 13974 23910 14026 23962
rect 16782 23910 16834 23962
rect 16846 23910 16898 23962
rect 16910 23910 16962 23962
rect 16974 23910 17026 23962
rect 19782 23910 19834 23962
rect 19846 23910 19898 23962
rect 19910 23910 19962 23962
rect 19974 23910 20026 23962
rect 22782 23910 22834 23962
rect 22846 23910 22898 23962
rect 22910 23910 22962 23962
rect 22974 23910 23026 23962
rect 25782 23910 25834 23962
rect 25846 23910 25898 23962
rect 25910 23910 25962 23962
rect 25974 23910 26026 23962
rect 3282 23366 3334 23418
rect 3346 23366 3398 23418
rect 3410 23366 3462 23418
rect 3474 23366 3526 23418
rect 6282 23366 6334 23418
rect 6346 23366 6398 23418
rect 6410 23366 6462 23418
rect 6474 23366 6526 23418
rect 9282 23366 9334 23418
rect 9346 23366 9398 23418
rect 9410 23366 9462 23418
rect 9474 23366 9526 23418
rect 12282 23366 12334 23418
rect 12346 23366 12398 23418
rect 12410 23366 12462 23418
rect 12474 23366 12526 23418
rect 15282 23366 15334 23418
rect 15346 23366 15398 23418
rect 15410 23366 15462 23418
rect 15474 23366 15526 23418
rect 18282 23366 18334 23418
rect 18346 23366 18398 23418
rect 18410 23366 18462 23418
rect 18474 23366 18526 23418
rect 21282 23366 21334 23418
rect 21346 23366 21398 23418
rect 21410 23366 21462 23418
rect 21474 23366 21526 23418
rect 24282 23366 24334 23418
rect 24346 23366 24398 23418
rect 24410 23366 24462 23418
rect 24474 23366 24526 23418
rect 27282 23366 27334 23418
rect 27346 23366 27398 23418
rect 27410 23366 27462 23418
rect 27474 23366 27526 23418
rect 1782 22822 1834 22874
rect 1846 22822 1898 22874
rect 1910 22822 1962 22874
rect 1974 22822 2026 22874
rect 4782 22822 4834 22874
rect 4846 22822 4898 22874
rect 4910 22822 4962 22874
rect 4974 22822 5026 22874
rect 7782 22822 7834 22874
rect 7846 22822 7898 22874
rect 7910 22822 7962 22874
rect 7974 22822 8026 22874
rect 10782 22822 10834 22874
rect 10846 22822 10898 22874
rect 10910 22822 10962 22874
rect 10974 22822 11026 22874
rect 13782 22822 13834 22874
rect 13846 22822 13898 22874
rect 13910 22822 13962 22874
rect 13974 22822 14026 22874
rect 16782 22822 16834 22874
rect 16846 22822 16898 22874
rect 16910 22822 16962 22874
rect 16974 22822 17026 22874
rect 19782 22822 19834 22874
rect 19846 22822 19898 22874
rect 19910 22822 19962 22874
rect 19974 22822 20026 22874
rect 22782 22822 22834 22874
rect 22846 22822 22898 22874
rect 22910 22822 22962 22874
rect 22974 22822 23026 22874
rect 25782 22822 25834 22874
rect 25846 22822 25898 22874
rect 25910 22822 25962 22874
rect 25974 22822 26026 22874
rect 3282 22278 3334 22330
rect 3346 22278 3398 22330
rect 3410 22278 3462 22330
rect 3474 22278 3526 22330
rect 6282 22278 6334 22330
rect 6346 22278 6398 22330
rect 6410 22278 6462 22330
rect 6474 22278 6526 22330
rect 9282 22278 9334 22330
rect 9346 22278 9398 22330
rect 9410 22278 9462 22330
rect 9474 22278 9526 22330
rect 12282 22278 12334 22330
rect 12346 22278 12398 22330
rect 12410 22278 12462 22330
rect 12474 22278 12526 22330
rect 15282 22278 15334 22330
rect 15346 22278 15398 22330
rect 15410 22278 15462 22330
rect 15474 22278 15526 22330
rect 18282 22278 18334 22330
rect 18346 22278 18398 22330
rect 18410 22278 18462 22330
rect 18474 22278 18526 22330
rect 21282 22278 21334 22330
rect 21346 22278 21398 22330
rect 21410 22278 21462 22330
rect 21474 22278 21526 22330
rect 24282 22278 24334 22330
rect 24346 22278 24398 22330
rect 24410 22278 24462 22330
rect 24474 22278 24526 22330
rect 27282 22278 27334 22330
rect 27346 22278 27398 22330
rect 27410 22278 27462 22330
rect 27474 22278 27526 22330
rect 1782 21734 1834 21786
rect 1846 21734 1898 21786
rect 1910 21734 1962 21786
rect 1974 21734 2026 21786
rect 4782 21734 4834 21786
rect 4846 21734 4898 21786
rect 4910 21734 4962 21786
rect 4974 21734 5026 21786
rect 7782 21734 7834 21786
rect 7846 21734 7898 21786
rect 7910 21734 7962 21786
rect 7974 21734 8026 21786
rect 10782 21734 10834 21786
rect 10846 21734 10898 21786
rect 10910 21734 10962 21786
rect 10974 21734 11026 21786
rect 13782 21734 13834 21786
rect 13846 21734 13898 21786
rect 13910 21734 13962 21786
rect 13974 21734 14026 21786
rect 16782 21734 16834 21786
rect 16846 21734 16898 21786
rect 16910 21734 16962 21786
rect 16974 21734 17026 21786
rect 19782 21734 19834 21786
rect 19846 21734 19898 21786
rect 19910 21734 19962 21786
rect 19974 21734 20026 21786
rect 22782 21734 22834 21786
rect 22846 21734 22898 21786
rect 22910 21734 22962 21786
rect 22974 21734 23026 21786
rect 25782 21734 25834 21786
rect 25846 21734 25898 21786
rect 25910 21734 25962 21786
rect 25974 21734 26026 21786
rect 3282 21190 3334 21242
rect 3346 21190 3398 21242
rect 3410 21190 3462 21242
rect 3474 21190 3526 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 6410 21190 6462 21242
rect 6474 21190 6526 21242
rect 9282 21190 9334 21242
rect 9346 21190 9398 21242
rect 9410 21190 9462 21242
rect 9474 21190 9526 21242
rect 12282 21190 12334 21242
rect 12346 21190 12398 21242
rect 12410 21190 12462 21242
rect 12474 21190 12526 21242
rect 15282 21190 15334 21242
rect 15346 21190 15398 21242
rect 15410 21190 15462 21242
rect 15474 21190 15526 21242
rect 18282 21190 18334 21242
rect 18346 21190 18398 21242
rect 18410 21190 18462 21242
rect 18474 21190 18526 21242
rect 21282 21190 21334 21242
rect 21346 21190 21398 21242
rect 21410 21190 21462 21242
rect 21474 21190 21526 21242
rect 24282 21190 24334 21242
rect 24346 21190 24398 21242
rect 24410 21190 24462 21242
rect 24474 21190 24526 21242
rect 27282 21190 27334 21242
rect 27346 21190 27398 21242
rect 27410 21190 27462 21242
rect 27474 21190 27526 21242
rect 1782 20646 1834 20698
rect 1846 20646 1898 20698
rect 1910 20646 1962 20698
rect 1974 20646 2026 20698
rect 4782 20646 4834 20698
rect 4846 20646 4898 20698
rect 4910 20646 4962 20698
rect 4974 20646 5026 20698
rect 7782 20646 7834 20698
rect 7846 20646 7898 20698
rect 7910 20646 7962 20698
rect 7974 20646 8026 20698
rect 10782 20646 10834 20698
rect 10846 20646 10898 20698
rect 10910 20646 10962 20698
rect 10974 20646 11026 20698
rect 13782 20646 13834 20698
rect 13846 20646 13898 20698
rect 13910 20646 13962 20698
rect 13974 20646 14026 20698
rect 16782 20646 16834 20698
rect 16846 20646 16898 20698
rect 16910 20646 16962 20698
rect 16974 20646 17026 20698
rect 19782 20646 19834 20698
rect 19846 20646 19898 20698
rect 19910 20646 19962 20698
rect 19974 20646 20026 20698
rect 22782 20646 22834 20698
rect 22846 20646 22898 20698
rect 22910 20646 22962 20698
rect 22974 20646 23026 20698
rect 25782 20646 25834 20698
rect 25846 20646 25898 20698
rect 25910 20646 25962 20698
rect 25974 20646 26026 20698
rect 3282 20102 3334 20154
rect 3346 20102 3398 20154
rect 3410 20102 3462 20154
rect 3474 20102 3526 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 6410 20102 6462 20154
rect 6474 20102 6526 20154
rect 9282 20102 9334 20154
rect 9346 20102 9398 20154
rect 9410 20102 9462 20154
rect 9474 20102 9526 20154
rect 12282 20102 12334 20154
rect 12346 20102 12398 20154
rect 12410 20102 12462 20154
rect 12474 20102 12526 20154
rect 15282 20102 15334 20154
rect 15346 20102 15398 20154
rect 15410 20102 15462 20154
rect 15474 20102 15526 20154
rect 18282 20102 18334 20154
rect 18346 20102 18398 20154
rect 18410 20102 18462 20154
rect 18474 20102 18526 20154
rect 21282 20102 21334 20154
rect 21346 20102 21398 20154
rect 21410 20102 21462 20154
rect 21474 20102 21526 20154
rect 24282 20102 24334 20154
rect 24346 20102 24398 20154
rect 24410 20102 24462 20154
rect 24474 20102 24526 20154
rect 27282 20102 27334 20154
rect 27346 20102 27398 20154
rect 27410 20102 27462 20154
rect 27474 20102 27526 20154
rect 1782 19558 1834 19610
rect 1846 19558 1898 19610
rect 1910 19558 1962 19610
rect 1974 19558 2026 19610
rect 4782 19558 4834 19610
rect 4846 19558 4898 19610
rect 4910 19558 4962 19610
rect 4974 19558 5026 19610
rect 7782 19558 7834 19610
rect 7846 19558 7898 19610
rect 7910 19558 7962 19610
rect 7974 19558 8026 19610
rect 10782 19558 10834 19610
rect 10846 19558 10898 19610
rect 10910 19558 10962 19610
rect 10974 19558 11026 19610
rect 13782 19558 13834 19610
rect 13846 19558 13898 19610
rect 13910 19558 13962 19610
rect 13974 19558 14026 19610
rect 16782 19558 16834 19610
rect 16846 19558 16898 19610
rect 16910 19558 16962 19610
rect 16974 19558 17026 19610
rect 19782 19558 19834 19610
rect 19846 19558 19898 19610
rect 19910 19558 19962 19610
rect 19974 19558 20026 19610
rect 22782 19558 22834 19610
rect 22846 19558 22898 19610
rect 22910 19558 22962 19610
rect 22974 19558 23026 19610
rect 25782 19558 25834 19610
rect 25846 19558 25898 19610
rect 25910 19558 25962 19610
rect 25974 19558 26026 19610
rect 3282 19014 3334 19066
rect 3346 19014 3398 19066
rect 3410 19014 3462 19066
rect 3474 19014 3526 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 6410 19014 6462 19066
rect 6474 19014 6526 19066
rect 9282 19014 9334 19066
rect 9346 19014 9398 19066
rect 9410 19014 9462 19066
rect 9474 19014 9526 19066
rect 12282 19014 12334 19066
rect 12346 19014 12398 19066
rect 12410 19014 12462 19066
rect 12474 19014 12526 19066
rect 15282 19014 15334 19066
rect 15346 19014 15398 19066
rect 15410 19014 15462 19066
rect 15474 19014 15526 19066
rect 18282 19014 18334 19066
rect 18346 19014 18398 19066
rect 18410 19014 18462 19066
rect 18474 19014 18526 19066
rect 21282 19014 21334 19066
rect 21346 19014 21398 19066
rect 21410 19014 21462 19066
rect 21474 19014 21526 19066
rect 24282 19014 24334 19066
rect 24346 19014 24398 19066
rect 24410 19014 24462 19066
rect 24474 19014 24526 19066
rect 27282 19014 27334 19066
rect 27346 19014 27398 19066
rect 27410 19014 27462 19066
rect 27474 19014 27526 19066
rect 1782 18470 1834 18522
rect 1846 18470 1898 18522
rect 1910 18470 1962 18522
rect 1974 18470 2026 18522
rect 4782 18470 4834 18522
rect 4846 18470 4898 18522
rect 4910 18470 4962 18522
rect 4974 18470 5026 18522
rect 7782 18470 7834 18522
rect 7846 18470 7898 18522
rect 7910 18470 7962 18522
rect 7974 18470 8026 18522
rect 10782 18470 10834 18522
rect 10846 18470 10898 18522
rect 10910 18470 10962 18522
rect 10974 18470 11026 18522
rect 13782 18470 13834 18522
rect 13846 18470 13898 18522
rect 13910 18470 13962 18522
rect 13974 18470 14026 18522
rect 16782 18470 16834 18522
rect 16846 18470 16898 18522
rect 16910 18470 16962 18522
rect 16974 18470 17026 18522
rect 19782 18470 19834 18522
rect 19846 18470 19898 18522
rect 19910 18470 19962 18522
rect 19974 18470 20026 18522
rect 22782 18470 22834 18522
rect 22846 18470 22898 18522
rect 22910 18470 22962 18522
rect 22974 18470 23026 18522
rect 25782 18470 25834 18522
rect 25846 18470 25898 18522
rect 25910 18470 25962 18522
rect 25974 18470 26026 18522
rect 3282 17926 3334 17978
rect 3346 17926 3398 17978
rect 3410 17926 3462 17978
rect 3474 17926 3526 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 6410 17926 6462 17978
rect 6474 17926 6526 17978
rect 9282 17926 9334 17978
rect 9346 17926 9398 17978
rect 9410 17926 9462 17978
rect 9474 17926 9526 17978
rect 12282 17926 12334 17978
rect 12346 17926 12398 17978
rect 12410 17926 12462 17978
rect 12474 17926 12526 17978
rect 15282 17926 15334 17978
rect 15346 17926 15398 17978
rect 15410 17926 15462 17978
rect 15474 17926 15526 17978
rect 18282 17926 18334 17978
rect 18346 17926 18398 17978
rect 18410 17926 18462 17978
rect 18474 17926 18526 17978
rect 21282 17926 21334 17978
rect 21346 17926 21398 17978
rect 21410 17926 21462 17978
rect 21474 17926 21526 17978
rect 24282 17926 24334 17978
rect 24346 17926 24398 17978
rect 24410 17926 24462 17978
rect 24474 17926 24526 17978
rect 27282 17926 27334 17978
rect 27346 17926 27398 17978
rect 27410 17926 27462 17978
rect 27474 17926 27526 17978
rect 1782 17382 1834 17434
rect 1846 17382 1898 17434
rect 1910 17382 1962 17434
rect 1974 17382 2026 17434
rect 4782 17382 4834 17434
rect 4846 17382 4898 17434
rect 4910 17382 4962 17434
rect 4974 17382 5026 17434
rect 7782 17382 7834 17434
rect 7846 17382 7898 17434
rect 7910 17382 7962 17434
rect 7974 17382 8026 17434
rect 10782 17382 10834 17434
rect 10846 17382 10898 17434
rect 10910 17382 10962 17434
rect 10974 17382 11026 17434
rect 13782 17382 13834 17434
rect 13846 17382 13898 17434
rect 13910 17382 13962 17434
rect 13974 17382 14026 17434
rect 16782 17382 16834 17434
rect 16846 17382 16898 17434
rect 16910 17382 16962 17434
rect 16974 17382 17026 17434
rect 19782 17382 19834 17434
rect 19846 17382 19898 17434
rect 19910 17382 19962 17434
rect 19974 17382 20026 17434
rect 22782 17382 22834 17434
rect 22846 17382 22898 17434
rect 22910 17382 22962 17434
rect 22974 17382 23026 17434
rect 25782 17382 25834 17434
rect 25846 17382 25898 17434
rect 25910 17382 25962 17434
rect 25974 17382 26026 17434
rect 3282 16838 3334 16890
rect 3346 16838 3398 16890
rect 3410 16838 3462 16890
rect 3474 16838 3526 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 6410 16838 6462 16890
rect 6474 16838 6526 16890
rect 9282 16838 9334 16890
rect 9346 16838 9398 16890
rect 9410 16838 9462 16890
rect 9474 16838 9526 16890
rect 12282 16838 12334 16890
rect 12346 16838 12398 16890
rect 12410 16838 12462 16890
rect 12474 16838 12526 16890
rect 15282 16838 15334 16890
rect 15346 16838 15398 16890
rect 15410 16838 15462 16890
rect 15474 16838 15526 16890
rect 18282 16838 18334 16890
rect 18346 16838 18398 16890
rect 18410 16838 18462 16890
rect 18474 16838 18526 16890
rect 21282 16838 21334 16890
rect 21346 16838 21398 16890
rect 21410 16838 21462 16890
rect 21474 16838 21526 16890
rect 24282 16838 24334 16890
rect 24346 16838 24398 16890
rect 24410 16838 24462 16890
rect 24474 16838 24526 16890
rect 27282 16838 27334 16890
rect 27346 16838 27398 16890
rect 27410 16838 27462 16890
rect 27474 16838 27526 16890
rect 14740 16668 14792 16720
rect 14280 16532 14332 16584
rect 16304 16532 16356 16584
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 17132 16532 17184 16584
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 16120 16396 16172 16448
rect 1782 16294 1834 16346
rect 1846 16294 1898 16346
rect 1910 16294 1962 16346
rect 1974 16294 2026 16346
rect 4782 16294 4834 16346
rect 4846 16294 4898 16346
rect 4910 16294 4962 16346
rect 4974 16294 5026 16346
rect 7782 16294 7834 16346
rect 7846 16294 7898 16346
rect 7910 16294 7962 16346
rect 7974 16294 8026 16346
rect 10782 16294 10834 16346
rect 10846 16294 10898 16346
rect 10910 16294 10962 16346
rect 10974 16294 11026 16346
rect 13782 16294 13834 16346
rect 13846 16294 13898 16346
rect 13910 16294 13962 16346
rect 13974 16294 14026 16346
rect 16782 16294 16834 16346
rect 16846 16294 16898 16346
rect 16910 16294 16962 16346
rect 16974 16294 17026 16346
rect 19782 16294 19834 16346
rect 19846 16294 19898 16346
rect 19910 16294 19962 16346
rect 19974 16294 20026 16346
rect 22782 16294 22834 16346
rect 22846 16294 22898 16346
rect 22910 16294 22962 16346
rect 22974 16294 23026 16346
rect 25782 16294 25834 16346
rect 25846 16294 25898 16346
rect 25910 16294 25962 16346
rect 25974 16294 26026 16346
rect 14372 16192 14424 16244
rect 14648 16124 14700 16176
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 16304 16192 16356 16244
rect 17960 16192 18012 16244
rect 14740 16124 14792 16133
rect 19892 16099 19944 16108
rect 19892 16065 19901 16099
rect 19901 16065 19935 16099
rect 19935 16065 19944 16099
rect 19892 16056 19944 16065
rect 16120 15988 16172 16040
rect 18144 15988 18196 16040
rect 19616 15988 19668 16040
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 17132 15895 17184 15904
rect 13820 15852 13872 15861
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 3282 15750 3334 15802
rect 3346 15750 3398 15802
rect 3410 15750 3462 15802
rect 3474 15750 3526 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 6410 15750 6462 15802
rect 6474 15750 6526 15802
rect 9282 15750 9334 15802
rect 9346 15750 9398 15802
rect 9410 15750 9462 15802
rect 9474 15750 9526 15802
rect 12282 15750 12334 15802
rect 12346 15750 12398 15802
rect 12410 15750 12462 15802
rect 12474 15750 12526 15802
rect 15282 15750 15334 15802
rect 15346 15750 15398 15802
rect 15410 15750 15462 15802
rect 15474 15750 15526 15802
rect 18282 15750 18334 15802
rect 18346 15750 18398 15802
rect 18410 15750 18462 15802
rect 18474 15750 18526 15802
rect 21282 15750 21334 15802
rect 21346 15750 21398 15802
rect 21410 15750 21462 15802
rect 21474 15750 21526 15802
rect 24282 15750 24334 15802
rect 24346 15750 24398 15802
rect 24410 15750 24462 15802
rect 24474 15750 24526 15802
rect 27282 15750 27334 15802
rect 27346 15750 27398 15802
rect 27410 15750 27462 15802
rect 27474 15750 27526 15802
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 13820 15512 13872 15564
rect 14280 15512 14332 15564
rect 17132 15512 17184 15564
rect 17408 15512 17460 15564
rect 19432 15512 19484 15564
rect 19892 15512 19944 15564
rect 20720 15512 20772 15564
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 14556 15444 14608 15496
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 17684 15444 17736 15496
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 18144 15444 18196 15453
rect 19156 15487 19208 15496
rect 19156 15453 19165 15487
rect 19165 15453 19199 15487
rect 19199 15453 19208 15487
rect 19156 15444 19208 15453
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 21272 15376 21324 15428
rect 21916 15376 21968 15428
rect 12992 15351 13044 15360
rect 12992 15317 13001 15351
rect 13001 15317 13035 15351
rect 13035 15317 13044 15351
rect 12992 15308 13044 15317
rect 13360 15308 13412 15360
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15936 15351 15988 15360
rect 15936 15317 15945 15351
rect 15945 15317 15979 15351
rect 15979 15317 15988 15351
rect 15936 15308 15988 15317
rect 19524 15308 19576 15360
rect 1782 15206 1834 15258
rect 1846 15206 1898 15258
rect 1910 15206 1962 15258
rect 1974 15206 2026 15258
rect 4782 15206 4834 15258
rect 4846 15206 4898 15258
rect 4910 15206 4962 15258
rect 4974 15206 5026 15258
rect 7782 15206 7834 15258
rect 7846 15206 7898 15258
rect 7910 15206 7962 15258
rect 7974 15206 8026 15258
rect 10782 15206 10834 15258
rect 10846 15206 10898 15258
rect 10910 15206 10962 15258
rect 10974 15206 11026 15258
rect 13782 15206 13834 15258
rect 13846 15206 13898 15258
rect 13910 15206 13962 15258
rect 13974 15206 14026 15258
rect 16782 15206 16834 15258
rect 16846 15206 16898 15258
rect 16910 15206 16962 15258
rect 16974 15206 17026 15258
rect 19782 15206 19834 15258
rect 19846 15206 19898 15258
rect 19910 15206 19962 15258
rect 19974 15206 20026 15258
rect 22782 15206 22834 15258
rect 22846 15206 22898 15258
rect 22910 15206 22962 15258
rect 22974 15206 23026 15258
rect 25782 15206 25834 15258
rect 25846 15206 25898 15258
rect 25910 15206 25962 15258
rect 25974 15206 26026 15258
rect 12808 15104 12860 15156
rect 14648 15104 14700 15156
rect 14740 15104 14792 15156
rect 21088 15104 21140 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 13360 15036 13412 15088
rect 18144 15036 18196 15088
rect 19156 15036 19208 15088
rect 20352 15036 20404 15088
rect 14188 14968 14240 15020
rect 15752 14968 15804 15020
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 17684 14900 17736 14952
rect 17960 14900 18012 14952
rect 17592 14832 17644 14884
rect 18972 14832 19024 14884
rect 20168 15011 20220 15020
rect 20168 14977 20177 15011
rect 20177 14977 20211 15011
rect 20211 14977 20220 15011
rect 20168 14968 20220 14977
rect 21640 14968 21692 15020
rect 21180 14900 21232 14952
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 17408 14764 17460 14816
rect 18880 14807 18932 14816
rect 18880 14773 18889 14807
rect 18889 14773 18923 14807
rect 18923 14773 18932 14807
rect 18880 14764 18932 14773
rect 3282 14662 3334 14714
rect 3346 14662 3398 14714
rect 3410 14662 3462 14714
rect 3474 14662 3526 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 6410 14662 6462 14714
rect 6474 14662 6526 14714
rect 9282 14662 9334 14714
rect 9346 14662 9398 14714
rect 9410 14662 9462 14714
rect 9474 14662 9526 14714
rect 12282 14662 12334 14714
rect 12346 14662 12398 14714
rect 12410 14662 12462 14714
rect 12474 14662 12526 14714
rect 15282 14662 15334 14714
rect 15346 14662 15398 14714
rect 15410 14662 15462 14714
rect 15474 14662 15526 14714
rect 18282 14662 18334 14714
rect 18346 14662 18398 14714
rect 18410 14662 18462 14714
rect 18474 14662 18526 14714
rect 21282 14662 21334 14714
rect 21346 14662 21398 14714
rect 21410 14662 21462 14714
rect 21474 14662 21526 14714
rect 24282 14662 24334 14714
rect 24346 14662 24398 14714
rect 24410 14662 24462 14714
rect 24474 14662 24526 14714
rect 27282 14662 27334 14714
rect 27346 14662 27398 14714
rect 27410 14662 27462 14714
rect 27474 14662 27526 14714
rect 14096 14560 14148 14612
rect 14556 14560 14608 14612
rect 17592 14560 17644 14612
rect 17960 14560 18012 14612
rect 20168 14560 20220 14612
rect 21180 14603 21232 14612
rect 21180 14569 21189 14603
rect 21189 14569 21223 14603
rect 21223 14569 21232 14603
rect 21180 14560 21232 14569
rect 21640 14560 21692 14612
rect 12900 14467 12952 14476
rect 12900 14433 12909 14467
rect 12909 14433 12943 14467
rect 12943 14433 12952 14467
rect 12900 14424 12952 14433
rect 14188 14467 14240 14476
rect 11520 14356 11572 14408
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 14372 14424 14424 14476
rect 15660 14424 15712 14476
rect 20260 14424 20312 14476
rect 21088 14424 21140 14476
rect 21916 14424 21968 14476
rect 23848 14424 23900 14476
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13544 14399 13596 14408
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 13636 14356 13688 14408
rect 15476 14399 15528 14408
rect 12716 14288 12768 14340
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 15936 14356 15988 14408
rect 16672 14356 16724 14408
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 18972 14356 19024 14408
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 19616 14356 19668 14408
rect 11428 14220 11480 14272
rect 12624 14220 12676 14272
rect 16396 14288 16448 14340
rect 20168 14356 20220 14408
rect 20536 14288 20588 14340
rect 22652 14331 22704 14340
rect 22652 14297 22661 14331
rect 22661 14297 22695 14331
rect 22695 14297 22704 14331
rect 22652 14288 22704 14297
rect 23112 14288 23164 14340
rect 17776 14220 17828 14272
rect 19064 14263 19116 14272
rect 19064 14229 19073 14263
rect 19073 14229 19107 14263
rect 19107 14229 19116 14263
rect 19064 14220 19116 14229
rect 19616 14220 19668 14272
rect 1782 14118 1834 14170
rect 1846 14118 1898 14170
rect 1910 14118 1962 14170
rect 1974 14118 2026 14170
rect 4782 14118 4834 14170
rect 4846 14118 4898 14170
rect 4910 14118 4962 14170
rect 4974 14118 5026 14170
rect 7782 14118 7834 14170
rect 7846 14118 7898 14170
rect 7910 14118 7962 14170
rect 7974 14118 8026 14170
rect 10782 14118 10834 14170
rect 10846 14118 10898 14170
rect 10910 14118 10962 14170
rect 10974 14118 11026 14170
rect 13782 14118 13834 14170
rect 13846 14118 13898 14170
rect 13910 14118 13962 14170
rect 13974 14118 14026 14170
rect 16782 14118 16834 14170
rect 16846 14118 16898 14170
rect 16910 14118 16962 14170
rect 16974 14118 17026 14170
rect 19782 14118 19834 14170
rect 19846 14118 19898 14170
rect 19910 14118 19962 14170
rect 19974 14118 20026 14170
rect 22782 14118 22834 14170
rect 22846 14118 22898 14170
rect 22910 14118 22962 14170
rect 22974 14118 23026 14170
rect 25782 14118 25834 14170
rect 25846 14118 25898 14170
rect 25910 14118 25962 14170
rect 25974 14118 26026 14170
rect 12992 14016 13044 14068
rect 13268 14016 13320 14068
rect 13636 14016 13688 14068
rect 15476 14016 15528 14068
rect 17316 14016 17368 14068
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 13360 13948 13412 14000
rect 15568 13991 15620 14000
rect 8484 13880 8536 13932
rect 13452 13880 13504 13932
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 15568 13957 15577 13991
rect 15577 13957 15611 13991
rect 15611 13957 15620 13991
rect 15568 13948 15620 13957
rect 15752 13880 15804 13932
rect 17592 13948 17644 14000
rect 19156 14016 19208 14068
rect 19432 14016 19484 14068
rect 18880 13880 18932 13932
rect 20352 14016 20404 14068
rect 23112 14059 23164 14068
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 20260 13948 20312 14000
rect 20996 13923 21048 13932
rect 13544 13812 13596 13864
rect 16120 13812 16172 13864
rect 16672 13812 16724 13864
rect 17408 13812 17460 13864
rect 19432 13812 19484 13864
rect 19616 13855 19668 13864
rect 19616 13821 19625 13855
rect 19625 13821 19659 13855
rect 19659 13821 19668 13855
rect 19616 13812 19668 13821
rect 20076 13744 20128 13796
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 20536 13855 20588 13864
rect 20536 13821 20545 13855
rect 20545 13821 20579 13855
rect 20579 13821 20588 13855
rect 20536 13812 20588 13821
rect 22100 13744 22152 13796
rect 8852 13676 8904 13728
rect 11520 13676 11572 13728
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 18696 13676 18748 13728
rect 20168 13676 20220 13728
rect 22652 13676 22704 13728
rect 3282 13574 3334 13626
rect 3346 13574 3398 13626
rect 3410 13574 3462 13626
rect 3474 13574 3526 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 6410 13574 6462 13626
rect 6474 13574 6526 13626
rect 9282 13574 9334 13626
rect 9346 13574 9398 13626
rect 9410 13574 9462 13626
rect 9474 13574 9526 13626
rect 12282 13574 12334 13626
rect 12346 13574 12398 13626
rect 12410 13574 12462 13626
rect 12474 13574 12526 13626
rect 15282 13574 15334 13626
rect 15346 13574 15398 13626
rect 15410 13574 15462 13626
rect 15474 13574 15526 13626
rect 18282 13574 18334 13626
rect 18346 13574 18398 13626
rect 18410 13574 18462 13626
rect 18474 13574 18526 13626
rect 21282 13574 21334 13626
rect 21346 13574 21398 13626
rect 21410 13574 21462 13626
rect 21474 13574 21526 13626
rect 24282 13574 24334 13626
rect 24346 13574 24398 13626
rect 24410 13574 24462 13626
rect 24474 13574 24526 13626
rect 27282 13574 27334 13626
rect 27346 13574 27398 13626
rect 27410 13574 27462 13626
rect 27474 13574 27526 13626
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 12716 13472 12768 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 18880 13472 18932 13524
rect 20260 13472 20312 13524
rect 20536 13515 20588 13524
rect 20536 13481 20545 13515
rect 20545 13481 20579 13515
rect 20579 13481 20588 13515
rect 20536 13472 20588 13481
rect 20996 13472 21048 13524
rect 14372 13404 14424 13456
rect 15568 13404 15620 13456
rect 19156 13404 19208 13456
rect 19432 13404 19484 13456
rect 13452 13379 13504 13388
rect 13452 13345 13461 13379
rect 13461 13345 13495 13379
rect 13495 13345 13504 13379
rect 13452 13336 13504 13345
rect 13636 13336 13688 13388
rect 14004 13336 14056 13388
rect 14188 13379 14240 13388
rect 14188 13345 14197 13379
rect 14197 13345 14231 13379
rect 14231 13345 14240 13379
rect 14188 13336 14240 13345
rect 16120 13336 16172 13388
rect 17224 13336 17276 13388
rect 14556 13268 14608 13320
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 19524 13268 19576 13320
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 14832 13200 14884 13252
rect 15108 13200 15160 13252
rect 17592 13243 17644 13252
rect 17592 13209 17601 13243
rect 17601 13209 17635 13243
rect 17635 13209 17644 13243
rect 17592 13200 17644 13209
rect 18788 13200 18840 13252
rect 8116 13132 8168 13184
rect 8484 13132 8536 13184
rect 11704 13132 11756 13184
rect 13544 13132 13596 13184
rect 20996 13132 21048 13184
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 1782 13030 1834 13082
rect 1846 13030 1898 13082
rect 1910 13030 1962 13082
rect 1974 13030 2026 13082
rect 4782 13030 4834 13082
rect 4846 13030 4898 13082
rect 4910 13030 4962 13082
rect 4974 13030 5026 13082
rect 7782 13030 7834 13082
rect 7846 13030 7898 13082
rect 7910 13030 7962 13082
rect 7974 13030 8026 13082
rect 10782 13030 10834 13082
rect 10846 13030 10898 13082
rect 10910 13030 10962 13082
rect 10974 13030 11026 13082
rect 13782 13030 13834 13082
rect 13846 13030 13898 13082
rect 13910 13030 13962 13082
rect 13974 13030 14026 13082
rect 16782 13030 16834 13082
rect 16846 13030 16898 13082
rect 16910 13030 16962 13082
rect 16974 13030 17026 13082
rect 19782 13030 19834 13082
rect 19846 13030 19898 13082
rect 19910 13030 19962 13082
rect 19974 13030 20026 13082
rect 22782 13030 22834 13082
rect 22846 13030 22898 13082
rect 22910 13030 22962 13082
rect 22974 13030 23026 13082
rect 25782 13030 25834 13082
rect 25846 13030 25898 13082
rect 25910 13030 25962 13082
rect 25974 13030 26026 13082
rect 11520 12928 11572 12980
rect 13268 12928 13320 12980
rect 9128 12835 9180 12844
rect 9128 12801 9137 12835
rect 9137 12801 9171 12835
rect 9171 12801 9180 12835
rect 9128 12792 9180 12801
rect 15568 12928 15620 12980
rect 17132 12928 17184 12980
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 19524 12971 19576 12980
rect 19524 12937 19533 12971
rect 19533 12937 19567 12971
rect 19567 12937 19576 12971
rect 19524 12928 19576 12937
rect 18604 12860 18656 12912
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 11796 12724 11848 12776
rect 13360 12724 13412 12776
rect 14188 12792 14240 12844
rect 16580 12835 16632 12844
rect 16580 12801 16589 12835
rect 16589 12801 16623 12835
rect 16623 12801 16632 12835
rect 16580 12792 16632 12801
rect 16764 12792 16816 12844
rect 17408 12792 17460 12844
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 16212 12724 16264 12776
rect 16672 12724 16724 12776
rect 18144 12724 18196 12776
rect 20628 12792 20680 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 22560 12792 22612 12844
rect 20260 12724 20312 12776
rect 22376 12767 22428 12776
rect 14280 12656 14332 12708
rect 13360 12588 13412 12640
rect 13452 12588 13504 12640
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 15844 12588 15896 12640
rect 17132 12588 17184 12640
rect 20168 12588 20220 12640
rect 22376 12733 22385 12767
rect 22385 12733 22419 12767
rect 22419 12733 22428 12767
rect 22376 12724 22428 12733
rect 23756 12656 23808 12708
rect 21088 12588 21140 12640
rect 23204 12631 23256 12640
rect 23204 12597 23213 12631
rect 23213 12597 23247 12631
rect 23247 12597 23256 12631
rect 23204 12588 23256 12597
rect 3282 12486 3334 12538
rect 3346 12486 3398 12538
rect 3410 12486 3462 12538
rect 3474 12486 3526 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 6410 12486 6462 12538
rect 6474 12486 6526 12538
rect 9282 12486 9334 12538
rect 9346 12486 9398 12538
rect 9410 12486 9462 12538
rect 9474 12486 9526 12538
rect 12282 12486 12334 12538
rect 12346 12486 12398 12538
rect 12410 12486 12462 12538
rect 12474 12486 12526 12538
rect 15282 12486 15334 12538
rect 15346 12486 15398 12538
rect 15410 12486 15462 12538
rect 15474 12486 15526 12538
rect 18282 12486 18334 12538
rect 18346 12486 18398 12538
rect 18410 12486 18462 12538
rect 18474 12486 18526 12538
rect 21282 12486 21334 12538
rect 21346 12486 21398 12538
rect 21410 12486 21462 12538
rect 21474 12486 21526 12538
rect 24282 12486 24334 12538
rect 24346 12486 24398 12538
rect 24410 12486 24462 12538
rect 24474 12486 24526 12538
rect 27282 12486 27334 12538
rect 27346 12486 27398 12538
rect 27410 12486 27462 12538
rect 27474 12486 27526 12538
rect 9128 12427 9180 12436
rect 9128 12393 9137 12427
rect 9137 12393 9171 12427
rect 9171 12393 9180 12427
rect 9128 12384 9180 12393
rect 11520 12384 11572 12436
rect 13636 12384 13688 12436
rect 14280 12427 14332 12436
rect 14280 12393 14289 12427
rect 14289 12393 14323 12427
rect 14323 12393 14332 12427
rect 14280 12384 14332 12393
rect 16672 12384 16724 12436
rect 17684 12427 17736 12436
rect 15936 12359 15988 12368
rect 15936 12325 15945 12359
rect 15945 12325 15979 12359
rect 15979 12325 15988 12359
rect 15936 12316 15988 12325
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 8668 12248 8720 12300
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 15844 12248 15896 12300
rect 17684 12393 17693 12427
rect 17693 12393 17727 12427
rect 17727 12393 17736 12427
rect 17684 12384 17736 12393
rect 17776 12384 17828 12436
rect 20260 12427 20312 12436
rect 20260 12393 20269 12427
rect 20269 12393 20303 12427
rect 20303 12393 20312 12427
rect 20260 12384 20312 12393
rect 23204 12384 23256 12436
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 11428 12180 11480 12232
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 17316 12180 17368 12232
rect 18604 12316 18656 12368
rect 18696 12316 18748 12368
rect 22652 12316 22704 12368
rect 28724 12316 28776 12368
rect 18880 12180 18932 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 22376 12223 22428 12232
rect 22376 12189 22385 12223
rect 22385 12189 22419 12223
rect 22419 12189 22428 12223
rect 22376 12180 22428 12189
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 22652 12180 22704 12232
rect 23756 12180 23808 12232
rect 9864 12112 9916 12164
rect 12256 12112 12308 12164
rect 12808 12044 12860 12096
rect 13728 12112 13780 12164
rect 18788 12155 18840 12164
rect 18788 12121 18797 12155
rect 18797 12121 18831 12155
rect 18831 12121 18840 12155
rect 18788 12112 18840 12121
rect 15108 12044 15160 12096
rect 20168 12044 20220 12096
rect 22008 12044 22060 12096
rect 1782 11942 1834 11994
rect 1846 11942 1898 11994
rect 1910 11942 1962 11994
rect 1974 11942 2026 11994
rect 4782 11942 4834 11994
rect 4846 11942 4898 11994
rect 4910 11942 4962 11994
rect 4974 11942 5026 11994
rect 7782 11942 7834 11994
rect 7846 11942 7898 11994
rect 7910 11942 7962 11994
rect 7974 11942 8026 11994
rect 10782 11942 10834 11994
rect 10846 11942 10898 11994
rect 10910 11942 10962 11994
rect 10974 11942 11026 11994
rect 13782 11942 13834 11994
rect 13846 11942 13898 11994
rect 13910 11942 13962 11994
rect 13974 11942 14026 11994
rect 16782 11942 16834 11994
rect 16846 11942 16898 11994
rect 16910 11942 16962 11994
rect 16974 11942 17026 11994
rect 19782 11942 19834 11994
rect 19846 11942 19898 11994
rect 19910 11942 19962 11994
rect 19974 11942 20026 11994
rect 22782 11942 22834 11994
rect 22846 11942 22898 11994
rect 22910 11942 22962 11994
rect 22974 11942 23026 11994
rect 25782 11942 25834 11994
rect 25846 11942 25898 11994
rect 25910 11942 25962 11994
rect 25974 11942 26026 11994
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 8300 11840 8352 11892
rect 12256 11840 12308 11892
rect 13268 11840 13320 11892
rect 13544 11840 13596 11892
rect 14556 11840 14608 11892
rect 16580 11883 16632 11892
rect 16580 11849 16589 11883
rect 16589 11849 16623 11883
rect 16623 11849 16632 11883
rect 16580 11840 16632 11849
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17316 11840 17368 11892
rect 18144 11840 18196 11892
rect 18788 11840 18840 11892
rect 22376 11840 22428 11892
rect 11796 11772 11848 11824
rect 14280 11772 14332 11824
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 9128 11636 9180 11688
rect 9588 11636 9640 11688
rect 11520 11704 11572 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 16488 11704 16540 11756
rect 17132 11704 17184 11756
rect 20720 11772 20772 11824
rect 20996 11815 21048 11824
rect 20996 11781 21005 11815
rect 21005 11781 21039 11815
rect 21039 11781 21048 11815
rect 20996 11772 21048 11781
rect 21088 11772 21140 11824
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 19708 11704 19760 11756
rect 20260 11704 20312 11756
rect 20444 11704 20496 11756
rect 22560 11704 22612 11756
rect 8576 11568 8628 11620
rect 14096 11636 14148 11688
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 18604 11636 18656 11688
rect 21088 11636 21140 11688
rect 11612 11568 11664 11620
rect 13176 11568 13228 11620
rect 11428 11500 11480 11552
rect 16304 11500 16356 11552
rect 16672 11500 16724 11552
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 20628 11500 20680 11552
rect 21824 11500 21876 11552
rect 22008 11543 22060 11552
rect 22008 11509 22017 11543
rect 22017 11509 22051 11543
rect 22051 11509 22060 11543
rect 22008 11500 22060 11509
rect 3282 11398 3334 11450
rect 3346 11398 3398 11450
rect 3410 11398 3462 11450
rect 3474 11398 3526 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 6410 11398 6462 11450
rect 6474 11398 6526 11450
rect 9282 11398 9334 11450
rect 9346 11398 9398 11450
rect 9410 11398 9462 11450
rect 9474 11398 9526 11450
rect 12282 11398 12334 11450
rect 12346 11398 12398 11450
rect 12410 11398 12462 11450
rect 12474 11398 12526 11450
rect 15282 11398 15334 11450
rect 15346 11398 15398 11450
rect 15410 11398 15462 11450
rect 15474 11398 15526 11450
rect 18282 11398 18334 11450
rect 18346 11398 18398 11450
rect 18410 11398 18462 11450
rect 18474 11398 18526 11450
rect 21282 11398 21334 11450
rect 21346 11398 21398 11450
rect 21410 11398 21462 11450
rect 21474 11398 21526 11450
rect 24282 11398 24334 11450
rect 24346 11398 24398 11450
rect 24410 11398 24462 11450
rect 24474 11398 24526 11450
rect 27282 11398 27334 11450
rect 27346 11398 27398 11450
rect 27410 11398 27462 11450
rect 27474 11398 27526 11450
rect 9772 11296 9824 11348
rect 12808 11296 12860 11348
rect 13176 11296 13228 11348
rect 9588 11228 9640 11280
rect 11336 11160 11388 11212
rect 13268 11160 13320 11212
rect 11612 11135 11664 11144
rect 11152 11024 11204 11076
rect 8576 10956 8628 11008
rect 10416 10999 10468 11008
rect 10416 10965 10425 10999
rect 10425 10965 10459 10999
rect 10459 10965 10468 10999
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 14924 11296 14976 11348
rect 16488 11296 16540 11348
rect 19708 11339 19760 11348
rect 13636 11228 13688 11280
rect 14280 11228 14332 11280
rect 14832 11271 14884 11280
rect 14832 11237 14841 11271
rect 14841 11237 14875 11271
rect 14875 11237 14884 11271
rect 14832 11228 14884 11237
rect 16212 11228 16264 11280
rect 14372 11160 14424 11212
rect 16028 11203 16080 11212
rect 16028 11169 16037 11203
rect 16037 11169 16071 11203
rect 16071 11169 16080 11203
rect 16028 11160 16080 11169
rect 16396 11160 16448 11212
rect 15660 11092 15712 11144
rect 15936 11092 15988 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 19708 11305 19717 11339
rect 19717 11305 19751 11339
rect 19751 11305 19760 11339
rect 19708 11296 19760 11305
rect 19984 11296 20036 11348
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 22652 11296 22704 11348
rect 21824 11228 21876 11280
rect 22468 11160 22520 11212
rect 15108 11024 15160 11076
rect 19248 11092 19300 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 10416 10956 10468 10965
rect 11888 10956 11940 11008
rect 11980 10956 12032 11008
rect 12624 10956 12676 11008
rect 14280 10956 14332 11008
rect 17132 10956 17184 11008
rect 19432 11024 19484 11076
rect 18604 10956 18656 11008
rect 21088 10999 21140 11008
rect 21088 10965 21097 10999
rect 21097 10965 21131 10999
rect 21131 10965 21140 10999
rect 21088 10956 21140 10965
rect 1782 10854 1834 10906
rect 1846 10854 1898 10906
rect 1910 10854 1962 10906
rect 1974 10854 2026 10906
rect 4782 10854 4834 10906
rect 4846 10854 4898 10906
rect 4910 10854 4962 10906
rect 4974 10854 5026 10906
rect 7782 10854 7834 10906
rect 7846 10854 7898 10906
rect 7910 10854 7962 10906
rect 7974 10854 8026 10906
rect 10782 10854 10834 10906
rect 10846 10854 10898 10906
rect 10910 10854 10962 10906
rect 10974 10854 11026 10906
rect 13782 10854 13834 10906
rect 13846 10854 13898 10906
rect 13910 10854 13962 10906
rect 13974 10854 14026 10906
rect 16782 10854 16834 10906
rect 16846 10854 16898 10906
rect 16910 10854 16962 10906
rect 16974 10854 17026 10906
rect 19782 10854 19834 10906
rect 19846 10854 19898 10906
rect 19910 10854 19962 10906
rect 19974 10854 20026 10906
rect 22782 10854 22834 10906
rect 22846 10854 22898 10906
rect 22910 10854 22962 10906
rect 22974 10854 23026 10906
rect 25782 10854 25834 10906
rect 25846 10854 25898 10906
rect 25910 10854 25962 10906
rect 25974 10854 26026 10906
rect 8300 10752 8352 10804
rect 8668 10684 8720 10736
rect 9036 10684 9088 10736
rect 8760 10659 8812 10668
rect 8760 10625 8769 10659
rect 8769 10625 8803 10659
rect 8803 10625 8812 10659
rect 8760 10616 8812 10625
rect 12164 10752 12216 10804
rect 16028 10795 16080 10804
rect 10324 10616 10376 10668
rect 8208 10548 8260 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 11336 10684 11388 10736
rect 11704 10684 11756 10736
rect 14464 10684 14516 10736
rect 16028 10761 16037 10795
rect 16037 10761 16071 10795
rect 16071 10761 16080 10795
rect 16028 10752 16080 10761
rect 16488 10684 16540 10736
rect 19432 10752 19484 10804
rect 19616 10795 19668 10804
rect 19616 10761 19625 10795
rect 19625 10761 19659 10795
rect 19659 10761 19668 10795
rect 19616 10752 19668 10761
rect 20720 10752 20772 10804
rect 21088 10684 21140 10736
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 15660 10616 15712 10668
rect 17592 10616 17644 10668
rect 19156 10616 19208 10668
rect 20444 10616 20496 10668
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 22468 10752 22520 10804
rect 13544 10548 13596 10600
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 20352 10548 20404 10600
rect 8576 10412 8628 10464
rect 8852 10412 8904 10464
rect 19248 10480 19300 10532
rect 21180 10480 21232 10532
rect 11612 10412 11664 10464
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 16764 10412 16816 10464
rect 17960 10412 18012 10464
rect 22008 10480 22060 10532
rect 21640 10455 21692 10464
rect 21640 10421 21649 10455
rect 21649 10421 21683 10455
rect 21683 10421 21692 10455
rect 21640 10412 21692 10421
rect 3282 10310 3334 10362
rect 3346 10310 3398 10362
rect 3410 10310 3462 10362
rect 3474 10310 3526 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 6410 10310 6462 10362
rect 6474 10310 6526 10362
rect 9282 10310 9334 10362
rect 9346 10310 9398 10362
rect 9410 10310 9462 10362
rect 9474 10310 9526 10362
rect 12282 10310 12334 10362
rect 12346 10310 12398 10362
rect 12410 10310 12462 10362
rect 12474 10310 12526 10362
rect 15282 10310 15334 10362
rect 15346 10310 15398 10362
rect 15410 10310 15462 10362
rect 15474 10310 15526 10362
rect 18282 10310 18334 10362
rect 18346 10310 18398 10362
rect 18410 10310 18462 10362
rect 18474 10310 18526 10362
rect 21282 10310 21334 10362
rect 21346 10310 21398 10362
rect 21410 10310 21462 10362
rect 21474 10310 21526 10362
rect 24282 10310 24334 10362
rect 24346 10310 24398 10362
rect 24410 10310 24462 10362
rect 24474 10310 24526 10362
rect 27282 10310 27334 10362
rect 27346 10310 27398 10362
rect 27410 10310 27462 10362
rect 27474 10310 27526 10362
rect 8760 10208 8812 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 14004 10208 14056 10260
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 20076 10208 20128 10260
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 20996 10208 21048 10260
rect 21180 10208 21232 10260
rect 9036 10183 9088 10192
rect 9036 10149 9045 10183
rect 9045 10149 9079 10183
rect 9079 10149 9088 10183
rect 9036 10140 9088 10149
rect 14464 10140 14516 10192
rect 16396 10140 16448 10192
rect 7104 10072 7156 10124
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 11520 10072 11572 10124
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 15660 10072 15712 10124
rect 7012 9979 7064 9988
rect 7012 9945 7021 9979
rect 7021 9945 7055 9979
rect 7055 9945 7064 9979
rect 7012 9936 7064 9945
rect 7472 9936 7524 9988
rect 8760 9979 8812 9988
rect 8760 9945 8769 9979
rect 8769 9945 8803 9979
rect 8803 9945 8812 9979
rect 8760 9936 8812 9945
rect 13636 10004 13688 10056
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 18972 10072 19024 10124
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 16764 10004 16816 10056
rect 17316 10047 17368 10056
rect 11428 9936 11480 9988
rect 11612 9936 11664 9988
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 19064 10004 19116 10056
rect 21916 10004 21968 10056
rect 18236 9979 18288 9988
rect 10600 9868 10652 9920
rect 18236 9945 18245 9979
rect 18245 9945 18279 9979
rect 18279 9945 18288 9979
rect 19248 9979 19300 9988
rect 18236 9936 18288 9945
rect 14188 9868 14240 9920
rect 17132 9868 17184 9920
rect 17408 9868 17460 9920
rect 18788 9868 18840 9920
rect 19248 9945 19257 9979
rect 19257 9945 19291 9979
rect 19291 9945 19300 9979
rect 19248 9936 19300 9945
rect 21732 9936 21784 9988
rect 22284 9979 22336 9988
rect 22284 9945 22293 9979
rect 22293 9945 22327 9979
rect 22327 9945 22336 9979
rect 22284 9936 22336 9945
rect 24032 9979 24084 9988
rect 19340 9868 19392 9920
rect 22652 9868 22704 9920
rect 24032 9945 24041 9979
rect 24041 9945 24075 9979
rect 24075 9945 24084 9979
rect 24032 9936 24084 9945
rect 1782 9766 1834 9818
rect 1846 9766 1898 9818
rect 1910 9766 1962 9818
rect 1974 9766 2026 9818
rect 4782 9766 4834 9818
rect 4846 9766 4898 9818
rect 4910 9766 4962 9818
rect 4974 9766 5026 9818
rect 7782 9766 7834 9818
rect 7846 9766 7898 9818
rect 7910 9766 7962 9818
rect 7974 9766 8026 9818
rect 10782 9766 10834 9818
rect 10846 9766 10898 9818
rect 10910 9766 10962 9818
rect 10974 9766 11026 9818
rect 13782 9766 13834 9818
rect 13846 9766 13898 9818
rect 13910 9766 13962 9818
rect 13974 9766 14026 9818
rect 16782 9766 16834 9818
rect 16846 9766 16898 9818
rect 16910 9766 16962 9818
rect 16974 9766 17026 9818
rect 19782 9766 19834 9818
rect 19846 9766 19898 9818
rect 19910 9766 19962 9818
rect 19974 9766 20026 9818
rect 22782 9766 22834 9818
rect 22846 9766 22898 9818
rect 22910 9766 22962 9818
rect 22974 9766 23026 9818
rect 25782 9766 25834 9818
rect 25846 9766 25898 9818
rect 25910 9766 25962 9818
rect 25974 9766 26026 9818
rect 7012 9664 7064 9716
rect 9864 9664 9916 9716
rect 11152 9664 11204 9716
rect 13636 9707 13688 9716
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 14096 9664 14148 9716
rect 14556 9664 14608 9716
rect 16212 9664 16264 9716
rect 17592 9707 17644 9716
rect 17592 9673 17601 9707
rect 17601 9673 17635 9707
rect 17635 9673 17644 9707
rect 17592 9664 17644 9673
rect 18236 9664 18288 9716
rect 11888 9596 11940 9648
rect 15660 9639 15712 9648
rect 15660 9605 15669 9639
rect 15669 9605 15703 9639
rect 15703 9605 15712 9639
rect 15660 9596 15712 9605
rect 18972 9596 19024 9648
rect 20812 9596 20864 9648
rect 22284 9664 22336 9716
rect 22652 9664 22704 9716
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 8576 9571 8628 9580
rect 8576 9537 8585 9571
rect 8585 9537 8619 9571
rect 8619 9537 8628 9571
rect 8576 9528 8628 9537
rect 9772 9528 9824 9580
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 10600 9528 10652 9580
rect 12900 9528 12952 9580
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 16304 9528 16356 9580
rect 9036 9503 9088 9512
rect 7472 9392 7524 9444
rect 9036 9469 9045 9503
rect 9045 9469 9079 9503
rect 9079 9469 9088 9503
rect 9036 9460 9088 9469
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 11704 9460 11756 9512
rect 16120 9460 16172 9512
rect 16580 9528 16632 9580
rect 19340 9571 19392 9580
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 19708 9571 19760 9580
rect 17316 9460 17368 9512
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 19524 9460 19576 9512
rect 20076 9528 20128 9580
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 21088 9528 21140 9580
rect 22652 9528 22704 9580
rect 24032 9528 24084 9580
rect 8760 9392 8812 9444
rect 11428 9435 11480 9444
rect 11428 9401 11437 9435
rect 11437 9401 11471 9435
rect 11471 9401 11480 9435
rect 11428 9392 11480 9401
rect 11888 9392 11940 9444
rect 13544 9392 13596 9444
rect 14188 9392 14240 9444
rect 16304 9392 16356 9444
rect 21180 9392 21232 9444
rect 22192 9392 22244 9444
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 9956 9324 10008 9376
rect 11612 9324 11664 9376
rect 16672 9324 16724 9376
rect 19064 9324 19116 9376
rect 21916 9324 21968 9376
rect 3282 9222 3334 9274
rect 3346 9222 3398 9274
rect 3410 9222 3462 9274
rect 3474 9222 3526 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 6410 9222 6462 9274
rect 6474 9222 6526 9274
rect 9282 9222 9334 9274
rect 9346 9222 9398 9274
rect 9410 9222 9462 9274
rect 9474 9222 9526 9274
rect 12282 9222 12334 9274
rect 12346 9222 12398 9274
rect 12410 9222 12462 9274
rect 12474 9222 12526 9274
rect 15282 9222 15334 9274
rect 15346 9222 15398 9274
rect 15410 9222 15462 9274
rect 15474 9222 15526 9274
rect 18282 9222 18334 9274
rect 18346 9222 18398 9274
rect 18410 9222 18462 9274
rect 18474 9222 18526 9274
rect 21282 9222 21334 9274
rect 21346 9222 21398 9274
rect 21410 9222 21462 9274
rect 21474 9222 21526 9274
rect 24282 9222 24334 9274
rect 24346 9222 24398 9274
rect 24410 9222 24462 9274
rect 24474 9222 24526 9274
rect 27282 9222 27334 9274
rect 27346 9222 27398 9274
rect 27410 9222 27462 9274
rect 27474 9222 27526 9274
rect 7472 9120 7524 9172
rect 8300 9120 8352 9172
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 11612 9120 11664 9172
rect 14280 9120 14332 9172
rect 14464 9163 14516 9172
rect 14464 9129 14473 9163
rect 14473 9129 14507 9163
rect 14507 9129 14516 9163
rect 14464 9120 14516 9129
rect 16212 9120 16264 9172
rect 19616 9120 19668 9172
rect 19708 9120 19760 9172
rect 22284 9163 22336 9172
rect 22284 9129 22293 9163
rect 22293 9129 22327 9163
rect 22327 9129 22336 9163
rect 22284 9120 22336 9129
rect 8208 9052 8260 9104
rect 10508 9052 10560 9104
rect 9128 8984 9180 9036
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10416 8984 10468 8993
rect 16028 8984 16080 9036
rect 16488 8984 16540 9036
rect 17408 9027 17460 9036
rect 17408 8993 17417 9027
rect 17417 8993 17451 9027
rect 17451 8993 17460 9027
rect 17408 8984 17460 8993
rect 19156 9027 19208 9036
rect 19156 8993 19165 9027
rect 19165 8993 19199 9027
rect 19199 8993 19208 9027
rect 19156 8984 19208 8993
rect 21088 9027 21140 9036
rect 21088 8993 21097 9027
rect 21097 8993 21131 9027
rect 21131 8993 21140 9027
rect 21088 8984 21140 8993
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 10324 8916 10376 8968
rect 11888 8916 11940 8968
rect 14372 8916 14424 8968
rect 15108 8916 15160 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 17132 8959 17184 8968
rect 15568 8916 15620 8925
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 21180 8916 21232 8968
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 22008 8959 22060 8968
rect 21824 8916 21876 8925
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 8576 8848 8628 8900
rect 9864 8891 9916 8900
rect 9864 8857 9873 8891
rect 9873 8857 9907 8891
rect 9907 8857 9916 8891
rect 9864 8848 9916 8857
rect 12716 8891 12768 8900
rect 12716 8857 12725 8891
rect 12725 8857 12759 8891
rect 12759 8857 12768 8891
rect 12716 8848 12768 8857
rect 16028 8891 16080 8900
rect 16028 8857 16037 8891
rect 16037 8857 16071 8891
rect 16071 8857 16080 8891
rect 16028 8848 16080 8857
rect 17868 8848 17920 8900
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 12900 8780 12952 8832
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 16580 8780 16632 8832
rect 20260 8780 20312 8832
rect 1782 8678 1834 8730
rect 1846 8678 1898 8730
rect 1910 8678 1962 8730
rect 1974 8678 2026 8730
rect 4782 8678 4834 8730
rect 4846 8678 4898 8730
rect 4910 8678 4962 8730
rect 4974 8678 5026 8730
rect 7782 8678 7834 8730
rect 7846 8678 7898 8730
rect 7910 8678 7962 8730
rect 7974 8678 8026 8730
rect 10782 8678 10834 8730
rect 10846 8678 10898 8730
rect 10910 8678 10962 8730
rect 10974 8678 11026 8730
rect 13782 8678 13834 8730
rect 13846 8678 13898 8730
rect 13910 8678 13962 8730
rect 13974 8678 14026 8730
rect 16782 8678 16834 8730
rect 16846 8678 16898 8730
rect 16910 8678 16962 8730
rect 16974 8678 17026 8730
rect 19782 8678 19834 8730
rect 19846 8678 19898 8730
rect 19910 8678 19962 8730
rect 19974 8678 20026 8730
rect 22782 8678 22834 8730
rect 22846 8678 22898 8730
rect 22910 8678 22962 8730
rect 22974 8678 23026 8730
rect 25782 8678 25834 8730
rect 25846 8678 25898 8730
rect 25910 8678 25962 8730
rect 25974 8678 26026 8730
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 9036 8508 9088 8560
rect 15568 8576 15620 8628
rect 17132 8576 17184 8628
rect 21180 8576 21232 8628
rect 22008 8576 22060 8628
rect 22652 8576 22704 8628
rect 12900 8508 12952 8560
rect 14924 8508 14976 8560
rect 8944 8440 8996 8492
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 10600 8440 10652 8492
rect 11704 8440 11756 8492
rect 12716 8440 12768 8492
rect 15108 8440 15160 8492
rect 16304 8440 16356 8492
rect 18144 8440 18196 8492
rect 20812 8508 20864 8560
rect 21640 8508 21692 8560
rect 19156 8440 19208 8492
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 19892 8483 19944 8492
rect 13268 8415 13320 8424
rect 5724 8236 5776 8288
rect 7196 8279 7248 8288
rect 7196 8245 7205 8279
rect 7205 8245 7239 8279
rect 7239 8245 7248 8279
rect 7196 8236 7248 8245
rect 7932 8279 7984 8288
rect 7932 8245 7941 8279
rect 7941 8245 7975 8279
rect 7975 8245 7984 8279
rect 7932 8236 7984 8245
rect 8300 8236 8352 8288
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 14464 8372 14516 8424
rect 19892 8449 19901 8483
rect 19901 8449 19935 8483
rect 19935 8449 19944 8483
rect 19892 8440 19944 8449
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20444 8483 20496 8492
rect 20444 8449 20462 8483
rect 20462 8449 20496 8483
rect 20444 8440 20496 8449
rect 21548 8440 21600 8492
rect 9864 8236 9916 8288
rect 11888 8236 11940 8288
rect 14004 8236 14056 8288
rect 15108 8236 15160 8288
rect 16304 8236 16356 8288
rect 17500 8236 17552 8288
rect 19064 8236 19116 8288
rect 20076 8372 20128 8424
rect 22468 8279 22520 8288
rect 22468 8245 22477 8279
rect 22477 8245 22511 8279
rect 22511 8245 22520 8279
rect 22468 8236 22520 8245
rect 3282 8134 3334 8186
rect 3346 8134 3398 8186
rect 3410 8134 3462 8186
rect 3474 8134 3526 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 6410 8134 6462 8186
rect 6474 8134 6526 8186
rect 9282 8134 9334 8186
rect 9346 8134 9398 8186
rect 9410 8134 9462 8186
rect 9474 8134 9526 8186
rect 12282 8134 12334 8186
rect 12346 8134 12398 8186
rect 12410 8134 12462 8186
rect 12474 8134 12526 8186
rect 15282 8134 15334 8186
rect 15346 8134 15398 8186
rect 15410 8134 15462 8186
rect 15474 8134 15526 8186
rect 18282 8134 18334 8186
rect 18346 8134 18398 8186
rect 18410 8134 18462 8186
rect 18474 8134 18526 8186
rect 21282 8134 21334 8186
rect 21346 8134 21398 8186
rect 21410 8134 21462 8186
rect 21474 8134 21526 8186
rect 24282 8134 24334 8186
rect 24346 8134 24398 8186
rect 24410 8134 24462 8186
rect 24474 8134 24526 8186
rect 27282 8134 27334 8186
rect 27346 8134 27398 8186
rect 27410 8134 27462 8186
rect 27474 8134 27526 8186
rect 8944 8032 8996 8084
rect 10048 8075 10100 8084
rect 10048 8041 10057 8075
rect 10057 8041 10091 8075
rect 10091 8041 10100 8075
rect 10048 8032 10100 8041
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 12716 8032 12768 8084
rect 14924 8075 14976 8084
rect 14924 8041 14933 8075
rect 14933 8041 14967 8075
rect 14967 8041 14976 8075
rect 14924 8032 14976 8041
rect 17408 8032 17460 8084
rect 18144 8032 18196 8084
rect 19064 8032 19116 8084
rect 19524 8032 19576 8084
rect 19616 8032 19668 8084
rect 21824 8032 21876 8084
rect 22468 8032 22520 8084
rect 7196 7964 7248 8016
rect 12900 7964 12952 8016
rect 18972 8007 19024 8016
rect 18972 7973 18981 8007
rect 18981 7973 19015 8007
rect 19015 7973 19024 8007
rect 18972 7964 19024 7973
rect 20260 7964 20312 8016
rect 6184 7896 6236 7948
rect 7932 7828 7984 7880
rect 9956 7896 10008 7948
rect 13268 7939 13320 7948
rect 13268 7905 13277 7939
rect 13277 7905 13311 7939
rect 13311 7905 13320 7939
rect 13268 7896 13320 7905
rect 7472 7760 7524 7812
rect 8944 7828 8996 7880
rect 8668 7760 8720 7812
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 15108 7896 15160 7948
rect 19616 7896 19668 7948
rect 21640 7896 21692 7948
rect 13820 7828 13872 7837
rect 14004 7828 14056 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 15844 7828 15896 7880
rect 16212 7828 16264 7880
rect 16672 7828 16724 7880
rect 18144 7828 18196 7880
rect 21732 7871 21784 7880
rect 17132 7803 17184 7812
rect 9864 7692 9916 7744
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 11244 7692 11296 7744
rect 17132 7769 17141 7803
rect 17141 7769 17175 7803
rect 17175 7769 17184 7803
rect 17132 7760 17184 7769
rect 17224 7760 17276 7812
rect 19892 7760 19944 7812
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 21824 7760 21876 7812
rect 15752 7692 15804 7744
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 18696 7692 18748 7744
rect 20444 7692 20496 7744
rect 1782 7590 1834 7642
rect 1846 7590 1898 7642
rect 1910 7590 1962 7642
rect 1974 7590 2026 7642
rect 4782 7590 4834 7642
rect 4846 7590 4898 7642
rect 4910 7590 4962 7642
rect 4974 7590 5026 7642
rect 7782 7590 7834 7642
rect 7846 7590 7898 7642
rect 7910 7590 7962 7642
rect 7974 7590 8026 7642
rect 10782 7590 10834 7642
rect 10846 7590 10898 7642
rect 10910 7590 10962 7642
rect 10974 7590 11026 7642
rect 13782 7590 13834 7642
rect 13846 7590 13898 7642
rect 13910 7590 13962 7642
rect 13974 7590 14026 7642
rect 16782 7590 16834 7642
rect 16846 7590 16898 7642
rect 16910 7590 16962 7642
rect 16974 7590 17026 7642
rect 19782 7590 19834 7642
rect 19846 7590 19898 7642
rect 19910 7590 19962 7642
rect 19974 7590 20026 7642
rect 22782 7590 22834 7642
rect 22846 7590 22898 7642
rect 22910 7590 22962 7642
rect 22974 7590 23026 7642
rect 25782 7590 25834 7642
rect 25846 7590 25898 7642
rect 25910 7590 25962 7642
rect 25974 7590 26026 7642
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 11244 7488 11296 7540
rect 13636 7488 13688 7540
rect 14280 7531 14332 7540
rect 14280 7497 14289 7531
rect 14289 7497 14323 7531
rect 14323 7497 14332 7531
rect 14280 7488 14332 7497
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 17224 7488 17276 7540
rect 18144 7488 18196 7540
rect 10048 7420 10100 7472
rect 15844 7420 15896 7472
rect 16396 7420 16448 7472
rect 19616 7488 19668 7540
rect 21732 7488 21784 7540
rect 21824 7463 21876 7472
rect 21824 7429 21833 7463
rect 21833 7429 21867 7463
rect 21867 7429 21876 7463
rect 21824 7420 21876 7429
rect 7472 7352 7524 7404
rect 9128 7352 9180 7404
rect 10324 7352 10376 7404
rect 11704 7352 11756 7404
rect 12900 7352 12952 7404
rect 13728 7352 13780 7404
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 17040 7352 17092 7404
rect 17500 7352 17552 7404
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 20996 7352 21048 7404
rect 21732 7352 21784 7404
rect 22284 7395 22336 7404
rect 22284 7361 22293 7395
rect 22293 7361 22327 7395
rect 22327 7361 22336 7395
rect 22284 7352 22336 7361
rect 9956 7284 10008 7336
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 20628 7284 20680 7336
rect 21180 7284 21232 7336
rect 13452 7216 13504 7268
rect 14280 7216 14332 7268
rect 7564 7148 7616 7200
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12072 7148 12124 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13084 7148 13136 7200
rect 15936 7148 15988 7200
rect 16672 7148 16724 7200
rect 20536 7191 20588 7200
rect 20536 7157 20545 7191
rect 20545 7157 20579 7191
rect 20579 7157 20588 7191
rect 20536 7148 20588 7157
rect 21180 7148 21232 7200
rect 21916 7148 21968 7200
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 3282 7046 3334 7098
rect 3346 7046 3398 7098
rect 3410 7046 3462 7098
rect 3474 7046 3526 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 6410 7046 6462 7098
rect 6474 7046 6526 7098
rect 9282 7046 9334 7098
rect 9346 7046 9398 7098
rect 9410 7046 9462 7098
rect 9474 7046 9526 7098
rect 12282 7046 12334 7098
rect 12346 7046 12398 7098
rect 12410 7046 12462 7098
rect 12474 7046 12526 7098
rect 15282 7046 15334 7098
rect 15346 7046 15398 7098
rect 15410 7046 15462 7098
rect 15474 7046 15526 7098
rect 18282 7046 18334 7098
rect 18346 7046 18398 7098
rect 18410 7046 18462 7098
rect 18474 7046 18526 7098
rect 21282 7046 21334 7098
rect 21346 7046 21398 7098
rect 21410 7046 21462 7098
rect 21474 7046 21526 7098
rect 24282 7046 24334 7098
rect 24346 7046 24398 7098
rect 24410 7046 24462 7098
rect 24474 7046 24526 7098
rect 27282 7046 27334 7098
rect 27346 7046 27398 7098
rect 27410 7046 27462 7098
rect 27474 7046 27526 7098
rect 13728 6944 13780 6996
rect 14188 6944 14240 6996
rect 17040 6987 17092 6996
rect 17040 6953 17049 6987
rect 17049 6953 17083 6987
rect 17083 6953 17092 6987
rect 17040 6944 17092 6953
rect 18972 6944 19024 6996
rect 20260 6944 20312 6996
rect 15568 6919 15620 6928
rect 15568 6885 15577 6919
rect 15577 6885 15611 6919
rect 15611 6885 15620 6919
rect 15568 6876 15620 6885
rect 15844 6876 15896 6928
rect 19064 6876 19116 6928
rect 7656 6808 7708 6860
rect 6736 6740 6788 6792
rect 7564 6740 7616 6792
rect 12624 6808 12676 6860
rect 13176 6808 13228 6860
rect 14280 6808 14332 6860
rect 16304 6808 16356 6860
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 19156 6808 19208 6860
rect 19524 6808 19576 6860
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8668 6783 8720 6792
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 10508 6783 10560 6792
rect 8668 6740 8720 6749
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11888 6740 11940 6792
rect 7380 6672 7432 6724
rect 9864 6672 9916 6724
rect 12624 6715 12676 6724
rect 12624 6681 12633 6715
rect 12633 6681 12667 6715
rect 12667 6681 12676 6715
rect 12624 6672 12676 6681
rect 13084 6672 13136 6724
rect 15936 6672 15988 6724
rect 18144 6740 18196 6792
rect 18604 6740 18656 6792
rect 19340 6740 19392 6792
rect 20076 6808 20128 6860
rect 20536 6808 20588 6860
rect 21088 6808 21140 6860
rect 21824 6808 21876 6860
rect 21180 6783 21232 6792
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 17592 6672 17644 6724
rect 21548 6672 21600 6724
rect 22468 6672 22520 6724
rect 7564 6604 7616 6656
rect 9128 6604 9180 6656
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 16488 6604 16540 6656
rect 18880 6604 18932 6656
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 1782 6502 1834 6554
rect 1846 6502 1898 6554
rect 1910 6502 1962 6554
rect 1974 6502 2026 6554
rect 4782 6502 4834 6554
rect 4846 6502 4898 6554
rect 4910 6502 4962 6554
rect 4974 6502 5026 6554
rect 7782 6502 7834 6554
rect 7846 6502 7898 6554
rect 7910 6502 7962 6554
rect 7974 6502 8026 6554
rect 10782 6502 10834 6554
rect 10846 6502 10898 6554
rect 10910 6502 10962 6554
rect 10974 6502 11026 6554
rect 13782 6502 13834 6554
rect 13846 6502 13898 6554
rect 13910 6502 13962 6554
rect 13974 6502 14026 6554
rect 16782 6502 16834 6554
rect 16846 6502 16898 6554
rect 16910 6502 16962 6554
rect 16974 6502 17026 6554
rect 19782 6502 19834 6554
rect 19846 6502 19898 6554
rect 19910 6502 19962 6554
rect 19974 6502 20026 6554
rect 22782 6502 22834 6554
rect 22846 6502 22898 6554
rect 22910 6502 22962 6554
rect 22974 6502 23026 6554
rect 25782 6502 25834 6554
rect 25846 6502 25898 6554
rect 25910 6502 25962 6554
rect 25974 6502 26026 6554
rect 7196 6400 7248 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 10508 6400 10560 6452
rect 13084 6400 13136 6452
rect 17592 6400 17644 6452
rect 20076 6400 20128 6452
rect 21548 6400 21600 6452
rect 22284 6400 22336 6452
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 8668 6264 8720 6316
rect 11336 6375 11388 6384
rect 11336 6341 11345 6375
rect 11345 6341 11379 6375
rect 11379 6341 11388 6375
rect 11336 6332 11388 6341
rect 12900 6332 12952 6384
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 14372 6264 14424 6316
rect 16028 6264 16080 6316
rect 17408 6332 17460 6384
rect 19064 6375 19116 6384
rect 19064 6341 19073 6375
rect 19073 6341 19107 6375
rect 19107 6341 19116 6375
rect 19064 6332 19116 6341
rect 19800 6332 19852 6384
rect 21640 6375 21692 6384
rect 21640 6341 21649 6375
rect 21649 6341 21683 6375
rect 21683 6341 21692 6375
rect 21640 6332 21692 6341
rect 16488 6264 16540 6316
rect 21732 6307 21784 6316
rect 21732 6273 21741 6307
rect 21741 6273 21775 6307
rect 21775 6273 21784 6307
rect 21732 6264 21784 6273
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 10508 6239 10560 6248
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 11152 6196 11204 6248
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 14280 6196 14332 6248
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 15936 6128 15988 6180
rect 18604 6196 18656 6248
rect 8116 6060 8168 6112
rect 11888 6060 11940 6112
rect 12992 6060 13044 6112
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 16120 6060 16172 6112
rect 18144 6060 18196 6112
rect 19156 6196 19208 6248
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 3282 5958 3334 6010
rect 3346 5958 3398 6010
rect 3410 5958 3462 6010
rect 3474 5958 3526 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 6410 5958 6462 6010
rect 6474 5958 6526 6010
rect 9282 5958 9334 6010
rect 9346 5958 9398 6010
rect 9410 5958 9462 6010
rect 9474 5958 9526 6010
rect 12282 5958 12334 6010
rect 12346 5958 12398 6010
rect 12410 5958 12462 6010
rect 12474 5958 12526 6010
rect 15282 5958 15334 6010
rect 15346 5958 15398 6010
rect 15410 5958 15462 6010
rect 15474 5958 15526 6010
rect 18282 5958 18334 6010
rect 18346 5958 18398 6010
rect 18410 5958 18462 6010
rect 18474 5958 18526 6010
rect 21282 5958 21334 6010
rect 21346 5958 21398 6010
rect 21410 5958 21462 6010
rect 21474 5958 21526 6010
rect 24282 5958 24334 6010
rect 24346 5958 24398 6010
rect 24410 5958 24462 6010
rect 24474 5958 24526 6010
rect 27282 5958 27334 6010
rect 27346 5958 27398 6010
rect 27410 5958 27462 6010
rect 27474 5958 27526 6010
rect 5724 5899 5776 5908
rect 5724 5865 5733 5899
rect 5733 5865 5767 5899
rect 5767 5865 5776 5899
rect 5724 5856 5776 5865
rect 6736 5856 6788 5908
rect 7380 5856 7432 5908
rect 7656 5856 7708 5908
rect 8576 5856 8628 5908
rect 12624 5856 12676 5908
rect 13084 5856 13136 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 19064 5856 19116 5908
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 20260 5856 20312 5908
rect 20996 5856 21048 5908
rect 21088 5856 21140 5908
rect 22468 5856 22520 5908
rect 9680 5788 9732 5840
rect 16028 5788 16080 5840
rect 10508 5720 10560 5772
rect 11980 5720 12032 5772
rect 13084 5720 13136 5772
rect 8116 5652 8168 5704
rect 9128 5652 9180 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 13176 5695 13228 5704
rect 12992 5652 13044 5661
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 18696 5720 18748 5772
rect 18880 5763 18932 5772
rect 18880 5729 18889 5763
rect 18889 5729 18923 5763
rect 18923 5729 18932 5763
rect 18880 5720 18932 5729
rect 20904 5720 20956 5772
rect 7656 5584 7708 5636
rect 9036 5584 9088 5636
rect 9864 5627 9916 5636
rect 9864 5593 9873 5627
rect 9873 5593 9907 5627
rect 9907 5593 9916 5627
rect 9864 5584 9916 5593
rect 11336 5584 11388 5636
rect 11796 5584 11848 5636
rect 14556 5652 14608 5704
rect 16672 5652 16724 5704
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 19156 5652 19208 5704
rect 15108 5584 15160 5636
rect 19248 5584 19300 5636
rect 7104 5516 7156 5568
rect 8852 5516 8904 5568
rect 14280 5516 14332 5568
rect 16028 5559 16080 5568
rect 16028 5525 16037 5559
rect 16037 5525 16071 5559
rect 16071 5525 16080 5559
rect 16028 5516 16080 5525
rect 16212 5516 16264 5568
rect 18604 5516 18656 5568
rect 21916 5559 21968 5568
rect 21916 5525 21925 5559
rect 21925 5525 21959 5559
rect 21959 5525 21968 5559
rect 21916 5516 21968 5525
rect 1782 5414 1834 5466
rect 1846 5414 1898 5466
rect 1910 5414 1962 5466
rect 1974 5414 2026 5466
rect 4782 5414 4834 5466
rect 4846 5414 4898 5466
rect 4910 5414 4962 5466
rect 4974 5414 5026 5466
rect 7782 5414 7834 5466
rect 7846 5414 7898 5466
rect 7910 5414 7962 5466
rect 7974 5414 8026 5466
rect 10782 5414 10834 5466
rect 10846 5414 10898 5466
rect 10910 5414 10962 5466
rect 10974 5414 11026 5466
rect 13782 5414 13834 5466
rect 13846 5414 13898 5466
rect 13910 5414 13962 5466
rect 13974 5414 14026 5466
rect 16782 5414 16834 5466
rect 16846 5414 16898 5466
rect 16910 5414 16962 5466
rect 16974 5414 17026 5466
rect 19782 5414 19834 5466
rect 19846 5414 19898 5466
rect 19910 5414 19962 5466
rect 19974 5414 20026 5466
rect 22782 5414 22834 5466
rect 22846 5414 22898 5466
rect 22910 5414 22962 5466
rect 22974 5414 23026 5466
rect 25782 5414 25834 5466
rect 25846 5414 25898 5466
rect 25910 5414 25962 5466
rect 25974 5414 26026 5466
rect 7196 5355 7248 5364
rect 7196 5321 7205 5355
rect 7205 5321 7239 5355
rect 7239 5321 7248 5355
rect 7196 5312 7248 5321
rect 7656 5312 7708 5364
rect 8668 5312 8720 5364
rect 9036 5355 9088 5364
rect 9036 5321 9045 5355
rect 9045 5321 9079 5355
rect 9079 5321 9088 5355
rect 9036 5312 9088 5321
rect 10048 5312 10100 5364
rect 10324 5312 10376 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 16488 5312 16540 5364
rect 16672 5312 16724 5364
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 20904 5355 20956 5364
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 21732 5355 21784 5364
rect 21732 5321 21741 5355
rect 21741 5321 21775 5355
rect 21775 5321 21784 5355
rect 21732 5312 21784 5321
rect 8944 5176 8996 5228
rect 9680 5176 9732 5228
rect 11428 5244 11480 5296
rect 16028 5244 16080 5296
rect 17592 5244 17644 5296
rect 18144 5244 18196 5296
rect 11152 5176 11204 5228
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 12072 5176 12124 5228
rect 14372 5176 14424 5228
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 17408 5176 17460 5228
rect 18604 5176 18656 5228
rect 20260 5287 20312 5296
rect 20260 5253 20269 5287
rect 20269 5253 20303 5287
rect 20303 5253 20312 5287
rect 20260 5244 20312 5253
rect 20168 5176 20220 5228
rect 11060 5108 11112 5160
rect 11520 5108 11572 5160
rect 11152 5040 11204 5092
rect 11704 5040 11756 5092
rect 12992 5108 13044 5160
rect 16304 5108 16356 5160
rect 17868 5108 17920 5160
rect 18696 5151 18748 5160
rect 18696 5117 18705 5151
rect 18705 5117 18739 5151
rect 18739 5117 18748 5151
rect 18696 5108 18748 5117
rect 19156 5108 19208 5160
rect 20444 5108 20496 5160
rect 21916 5108 21968 5160
rect 8760 4972 8812 5024
rect 9680 4972 9732 5024
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 16396 4972 16448 5024
rect 3282 4870 3334 4922
rect 3346 4870 3398 4922
rect 3410 4870 3462 4922
rect 3474 4870 3526 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 6410 4870 6462 4922
rect 6474 4870 6526 4922
rect 9282 4870 9334 4922
rect 9346 4870 9398 4922
rect 9410 4870 9462 4922
rect 9474 4870 9526 4922
rect 12282 4870 12334 4922
rect 12346 4870 12398 4922
rect 12410 4870 12462 4922
rect 12474 4870 12526 4922
rect 15282 4870 15334 4922
rect 15346 4870 15398 4922
rect 15410 4870 15462 4922
rect 15474 4870 15526 4922
rect 18282 4870 18334 4922
rect 18346 4870 18398 4922
rect 18410 4870 18462 4922
rect 18474 4870 18526 4922
rect 21282 4870 21334 4922
rect 21346 4870 21398 4922
rect 21410 4870 21462 4922
rect 21474 4870 21526 4922
rect 24282 4870 24334 4922
rect 24346 4870 24398 4922
rect 24410 4870 24462 4922
rect 24474 4870 24526 4922
rect 27282 4870 27334 4922
rect 27346 4870 27398 4922
rect 27410 4870 27462 4922
rect 27474 4870 27526 4922
rect 8116 4768 8168 4820
rect 11060 4768 11112 4820
rect 13636 4768 13688 4820
rect 14556 4811 14608 4820
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 18144 4811 18196 4820
rect 14556 4768 14608 4777
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 18880 4768 18932 4820
rect 19616 4768 19668 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 11336 4700 11388 4752
rect 15384 4700 15436 4752
rect 8208 4675 8260 4684
rect 8208 4641 8217 4675
rect 8217 4641 8251 4675
rect 8251 4641 8260 4675
rect 8208 4632 8260 4641
rect 11428 4632 11480 4684
rect 15108 4632 15160 4684
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 10416 4496 10468 4548
rect 11612 4564 11664 4616
rect 14188 4564 14240 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 17224 4564 17276 4616
rect 18144 4564 18196 4616
rect 18604 4564 18656 4616
rect 19616 4564 19668 4616
rect 11888 4496 11940 4548
rect 8944 4428 8996 4480
rect 11980 4428 12032 4480
rect 14372 4428 14424 4480
rect 16396 4496 16448 4548
rect 18788 4496 18840 4548
rect 1782 4326 1834 4378
rect 1846 4326 1898 4378
rect 1910 4326 1962 4378
rect 1974 4326 2026 4378
rect 4782 4326 4834 4378
rect 4846 4326 4898 4378
rect 4910 4326 4962 4378
rect 4974 4326 5026 4378
rect 7782 4326 7834 4378
rect 7846 4326 7898 4378
rect 7910 4326 7962 4378
rect 7974 4326 8026 4378
rect 10782 4326 10834 4378
rect 10846 4326 10898 4378
rect 10910 4326 10962 4378
rect 10974 4326 11026 4378
rect 13782 4326 13834 4378
rect 13846 4326 13898 4378
rect 13910 4326 13962 4378
rect 13974 4326 14026 4378
rect 16782 4326 16834 4378
rect 16846 4326 16898 4378
rect 16910 4326 16962 4378
rect 16974 4326 17026 4378
rect 19782 4326 19834 4378
rect 19846 4326 19898 4378
rect 19910 4326 19962 4378
rect 19974 4326 20026 4378
rect 22782 4326 22834 4378
rect 22846 4326 22898 4378
rect 22910 4326 22962 4378
rect 22974 4326 23026 4378
rect 25782 4326 25834 4378
rect 25846 4326 25898 4378
rect 25910 4326 25962 4378
rect 25974 4326 26026 4378
rect 8208 4224 8260 4276
rect 12624 4224 12676 4276
rect 14096 4224 14148 4276
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 19524 4224 19576 4276
rect 20444 4267 20496 4276
rect 20444 4233 20453 4267
rect 20453 4233 20487 4267
rect 20487 4233 20496 4267
rect 20444 4224 20496 4233
rect 9680 4156 9732 4208
rect 11244 4156 11296 4208
rect 11612 4156 11664 4208
rect 13544 4156 13596 4208
rect 14464 4156 14516 4208
rect 16672 4156 16724 4208
rect 8116 4131 8168 4140
rect 8116 4097 8125 4131
rect 8125 4097 8159 4131
rect 8159 4097 8168 4131
rect 8116 4088 8168 4097
rect 8760 4088 8812 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 15384 4131 15436 4140
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 8852 4020 8904 4072
rect 9128 4020 9180 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10140 4020 10192 4072
rect 11244 4020 11296 4072
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 18144 4088 18196 4140
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 19616 4131 19668 4140
rect 19616 4097 19625 4131
rect 19625 4097 19659 4131
rect 19659 4097 19668 4131
rect 19616 4088 19668 4097
rect 14096 4020 14148 4072
rect 11244 3884 11296 3936
rect 13176 3884 13228 3936
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 17224 3952 17276 4004
rect 15016 3884 15068 3936
rect 15844 3884 15896 3936
rect 16212 3884 16264 3936
rect 3282 3782 3334 3834
rect 3346 3782 3398 3834
rect 3410 3782 3462 3834
rect 3474 3782 3526 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 6410 3782 6462 3834
rect 6474 3782 6526 3834
rect 9282 3782 9334 3834
rect 9346 3782 9398 3834
rect 9410 3782 9462 3834
rect 9474 3782 9526 3834
rect 12282 3782 12334 3834
rect 12346 3782 12398 3834
rect 12410 3782 12462 3834
rect 12474 3782 12526 3834
rect 15282 3782 15334 3834
rect 15346 3782 15398 3834
rect 15410 3782 15462 3834
rect 15474 3782 15526 3834
rect 18282 3782 18334 3834
rect 18346 3782 18398 3834
rect 18410 3782 18462 3834
rect 18474 3782 18526 3834
rect 21282 3782 21334 3834
rect 21346 3782 21398 3834
rect 21410 3782 21462 3834
rect 21474 3782 21526 3834
rect 24282 3782 24334 3834
rect 24346 3782 24398 3834
rect 24410 3782 24462 3834
rect 24474 3782 24526 3834
rect 27282 3782 27334 3834
rect 27346 3782 27398 3834
rect 27410 3782 27462 3834
rect 27474 3782 27526 3834
rect 8760 3680 8812 3732
rect 8116 3612 8168 3664
rect 10232 3680 10284 3732
rect 11888 3680 11940 3732
rect 13636 3680 13688 3732
rect 16120 3680 16172 3732
rect 18696 3680 18748 3732
rect 15568 3655 15620 3664
rect 15568 3621 15577 3655
rect 15577 3621 15611 3655
rect 15611 3621 15620 3655
rect 15568 3612 15620 3621
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 17224 3544 17276 3596
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 19064 3544 19116 3596
rect 13636 3519 13688 3528
rect 9772 3408 9824 3460
rect 9128 3340 9180 3392
rect 10416 3451 10468 3460
rect 10416 3417 10425 3451
rect 10425 3417 10459 3451
rect 10459 3417 10468 3451
rect 10416 3408 10468 3417
rect 10508 3408 10560 3460
rect 12164 3451 12216 3460
rect 12164 3417 12173 3451
rect 12173 3417 12207 3451
rect 12207 3417 12216 3451
rect 12164 3408 12216 3417
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 16212 3476 16264 3528
rect 18604 3476 18656 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 16304 3408 16356 3460
rect 17776 3408 17828 3460
rect 13176 3383 13228 3392
rect 13176 3349 13185 3383
rect 13185 3349 13219 3383
rect 13219 3349 13228 3383
rect 13176 3340 13228 3349
rect 15016 3340 15068 3392
rect 1782 3238 1834 3290
rect 1846 3238 1898 3290
rect 1910 3238 1962 3290
rect 1974 3238 2026 3290
rect 4782 3238 4834 3290
rect 4846 3238 4898 3290
rect 4910 3238 4962 3290
rect 4974 3238 5026 3290
rect 7782 3238 7834 3290
rect 7846 3238 7898 3290
rect 7910 3238 7962 3290
rect 7974 3238 8026 3290
rect 10782 3238 10834 3290
rect 10846 3238 10898 3290
rect 10910 3238 10962 3290
rect 10974 3238 11026 3290
rect 13782 3238 13834 3290
rect 13846 3238 13898 3290
rect 13910 3238 13962 3290
rect 13974 3238 14026 3290
rect 16782 3238 16834 3290
rect 16846 3238 16898 3290
rect 16910 3238 16962 3290
rect 16974 3238 17026 3290
rect 19782 3238 19834 3290
rect 19846 3238 19898 3290
rect 19910 3238 19962 3290
rect 19974 3238 20026 3290
rect 22782 3238 22834 3290
rect 22846 3238 22898 3290
rect 22910 3238 22962 3290
rect 22974 3238 23026 3290
rect 25782 3238 25834 3290
rect 25846 3238 25898 3290
rect 25910 3238 25962 3290
rect 25974 3238 26026 3290
rect 8760 3136 8812 3188
rect 12072 3136 12124 3188
rect 17224 3136 17276 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 9772 3111 9824 3120
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 10232 3068 10284 3120
rect 8668 3000 8720 3052
rect 10140 3000 10192 3052
rect 13176 3068 13228 3120
rect 14464 3068 14516 3120
rect 11336 3000 11388 3052
rect 12624 3043 12676 3052
rect 12624 3009 12633 3043
rect 12633 3009 12667 3043
rect 12667 3009 12676 3043
rect 12624 3000 12676 3009
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 18144 3000 18196 3052
rect 10968 2932 11020 2984
rect 13728 2975 13780 2984
rect 10784 2864 10836 2916
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 14096 2932 14148 2984
rect 15016 2932 15068 2984
rect 15568 2864 15620 2916
rect 18604 2864 18656 2916
rect 10508 2796 10560 2848
rect 13728 2796 13780 2848
rect 16212 2839 16264 2848
rect 16212 2805 16221 2839
rect 16221 2805 16255 2839
rect 16255 2805 16264 2839
rect 16212 2796 16264 2805
rect 16304 2796 16356 2848
rect 3282 2694 3334 2746
rect 3346 2694 3398 2746
rect 3410 2694 3462 2746
rect 3474 2694 3526 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 6410 2694 6462 2746
rect 6474 2694 6526 2746
rect 9282 2694 9334 2746
rect 9346 2694 9398 2746
rect 9410 2694 9462 2746
rect 9474 2694 9526 2746
rect 12282 2694 12334 2746
rect 12346 2694 12398 2746
rect 12410 2694 12462 2746
rect 12474 2694 12526 2746
rect 15282 2694 15334 2746
rect 15346 2694 15398 2746
rect 15410 2694 15462 2746
rect 15474 2694 15526 2746
rect 18282 2694 18334 2746
rect 18346 2694 18398 2746
rect 18410 2694 18462 2746
rect 18474 2694 18526 2746
rect 21282 2694 21334 2746
rect 21346 2694 21398 2746
rect 21410 2694 21462 2746
rect 21474 2694 21526 2746
rect 24282 2694 24334 2746
rect 24346 2694 24398 2746
rect 24410 2694 24462 2746
rect 24474 2694 24526 2746
rect 27282 2694 27334 2746
rect 27346 2694 27398 2746
rect 27410 2694 27462 2746
rect 27474 2694 27526 2746
rect 8668 2592 8720 2644
rect 10508 2592 10560 2644
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 14464 2592 14516 2644
rect 17776 2592 17828 2644
rect 10416 2567 10468 2576
rect 10416 2533 10425 2567
rect 10425 2533 10459 2567
rect 10459 2533 10468 2567
rect 10416 2524 10468 2533
rect 13544 2524 13596 2576
rect 11152 2456 11204 2508
rect 11336 2456 11388 2508
rect 12164 2456 12216 2508
rect 15016 2456 15068 2508
rect 16672 2456 16724 2508
rect 18696 2456 18748 2508
rect 8944 2388 8996 2440
rect 10784 2388 10836 2440
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 11244 2431 11296 2440
rect 11244 2397 11253 2431
rect 11253 2397 11287 2431
rect 11287 2397 11296 2431
rect 11244 2388 11296 2397
rect 12072 2388 12124 2440
rect 13728 2388 13780 2440
rect 18236 2388 18288 2440
rect 18604 2388 18656 2440
rect 11244 2252 11296 2304
rect 14372 2320 14424 2372
rect 18144 2320 18196 2372
rect 14188 2252 14240 2304
rect 1782 2150 1834 2202
rect 1846 2150 1898 2202
rect 1910 2150 1962 2202
rect 1974 2150 2026 2202
rect 4782 2150 4834 2202
rect 4846 2150 4898 2202
rect 4910 2150 4962 2202
rect 4974 2150 5026 2202
rect 7782 2150 7834 2202
rect 7846 2150 7898 2202
rect 7910 2150 7962 2202
rect 7974 2150 8026 2202
rect 10782 2150 10834 2202
rect 10846 2150 10898 2202
rect 10910 2150 10962 2202
rect 10974 2150 11026 2202
rect 13782 2150 13834 2202
rect 13846 2150 13898 2202
rect 13910 2150 13962 2202
rect 13974 2150 14026 2202
rect 16782 2150 16834 2202
rect 16846 2150 16898 2202
rect 16910 2150 16962 2202
rect 16974 2150 17026 2202
rect 19782 2150 19834 2202
rect 19846 2150 19898 2202
rect 19910 2150 19962 2202
rect 19974 2150 20026 2202
rect 22782 2150 22834 2202
rect 22846 2150 22898 2202
rect 22910 2150 22962 2202
rect 22974 2150 23026 2202
rect 25782 2150 25834 2202
rect 25846 2150 25898 2202
rect 25910 2150 25962 2202
rect 25974 2150 26026 2202
rect 296 1300 348 1352
rect 10324 1300 10376 1352
<< metal2 >>
rect 6366 30871 6422 31671
rect 15658 30871 15714 31671
rect 24858 30954 24914 31671
rect 24596 30926 24914 30954
rect 1756 29404 2052 29424
rect 1812 29402 1836 29404
rect 1892 29402 1916 29404
rect 1972 29402 1996 29404
rect 1834 29350 1836 29402
rect 1898 29350 1910 29402
rect 1972 29350 1974 29402
rect 1812 29348 1836 29350
rect 1892 29348 1916 29350
rect 1972 29348 1996 29350
rect 1756 29328 2052 29348
rect 4756 29404 5052 29424
rect 4812 29402 4836 29404
rect 4892 29402 4916 29404
rect 4972 29402 4996 29404
rect 4834 29350 4836 29402
rect 4898 29350 4910 29402
rect 4972 29350 4974 29402
rect 4812 29348 4836 29350
rect 4892 29348 4916 29350
rect 4972 29348 4996 29350
rect 4756 29328 5052 29348
rect 7756 29404 8052 29424
rect 7812 29402 7836 29404
rect 7892 29402 7916 29404
rect 7972 29402 7996 29404
rect 7834 29350 7836 29402
rect 7898 29350 7910 29402
rect 7972 29350 7974 29402
rect 7812 29348 7836 29350
rect 7892 29348 7916 29350
rect 7972 29348 7996 29350
rect 7756 29328 8052 29348
rect 10756 29404 11052 29424
rect 10812 29402 10836 29404
rect 10892 29402 10916 29404
rect 10972 29402 10996 29404
rect 10834 29350 10836 29402
rect 10898 29350 10910 29402
rect 10972 29350 10974 29402
rect 10812 29348 10836 29350
rect 10892 29348 10916 29350
rect 10972 29348 10996 29350
rect 10756 29328 11052 29348
rect 13756 29404 14052 29424
rect 13812 29402 13836 29404
rect 13892 29402 13916 29404
rect 13972 29402 13996 29404
rect 13834 29350 13836 29402
rect 13898 29350 13910 29402
rect 13972 29350 13974 29402
rect 13812 29348 13836 29350
rect 13892 29348 13916 29350
rect 13972 29348 13996 29350
rect 13756 29328 14052 29348
rect 16756 29404 17052 29424
rect 16812 29402 16836 29404
rect 16892 29402 16916 29404
rect 16972 29402 16996 29404
rect 16834 29350 16836 29402
rect 16898 29350 16910 29402
rect 16972 29350 16974 29402
rect 16812 29348 16836 29350
rect 16892 29348 16916 29350
rect 16972 29348 16996 29350
rect 16756 29328 17052 29348
rect 19756 29404 20052 29424
rect 19812 29402 19836 29404
rect 19892 29402 19916 29404
rect 19972 29402 19996 29404
rect 19834 29350 19836 29402
rect 19898 29350 19910 29402
rect 19972 29350 19974 29402
rect 19812 29348 19836 29350
rect 19892 29348 19916 29350
rect 19972 29348 19996 29350
rect 19756 29328 20052 29348
rect 22756 29404 23052 29424
rect 22812 29402 22836 29404
rect 22892 29402 22916 29404
rect 22972 29402 22996 29404
rect 22834 29350 22836 29402
rect 22898 29350 22910 29402
rect 22972 29350 22974 29402
rect 22812 29348 22836 29350
rect 22892 29348 22916 29350
rect 22972 29348 22996 29350
rect 22756 29328 23052 29348
rect 3256 28860 3552 28880
rect 3312 28858 3336 28860
rect 3392 28858 3416 28860
rect 3472 28858 3496 28860
rect 3334 28806 3336 28858
rect 3398 28806 3410 28858
rect 3472 28806 3474 28858
rect 3312 28804 3336 28806
rect 3392 28804 3416 28806
rect 3472 28804 3496 28806
rect 3256 28784 3552 28804
rect 6256 28860 6552 28880
rect 6312 28858 6336 28860
rect 6392 28858 6416 28860
rect 6472 28858 6496 28860
rect 6334 28806 6336 28858
rect 6398 28806 6410 28858
rect 6472 28806 6474 28858
rect 6312 28804 6336 28806
rect 6392 28804 6416 28806
rect 6472 28804 6496 28806
rect 6256 28784 6552 28804
rect 9256 28860 9552 28880
rect 9312 28858 9336 28860
rect 9392 28858 9416 28860
rect 9472 28858 9496 28860
rect 9334 28806 9336 28858
rect 9398 28806 9410 28858
rect 9472 28806 9474 28858
rect 9312 28804 9336 28806
rect 9392 28804 9416 28806
rect 9472 28804 9496 28806
rect 9256 28784 9552 28804
rect 12256 28860 12552 28880
rect 12312 28858 12336 28860
rect 12392 28858 12416 28860
rect 12472 28858 12496 28860
rect 12334 28806 12336 28858
rect 12398 28806 12410 28858
rect 12472 28806 12474 28858
rect 12312 28804 12336 28806
rect 12392 28804 12416 28806
rect 12472 28804 12496 28806
rect 12256 28784 12552 28804
rect 15256 28860 15552 28880
rect 15312 28858 15336 28860
rect 15392 28858 15416 28860
rect 15472 28858 15496 28860
rect 15334 28806 15336 28858
rect 15398 28806 15410 28858
rect 15472 28806 15474 28858
rect 15312 28804 15336 28806
rect 15392 28804 15416 28806
rect 15472 28804 15496 28806
rect 15256 28784 15552 28804
rect 18256 28860 18552 28880
rect 18312 28858 18336 28860
rect 18392 28858 18416 28860
rect 18472 28858 18496 28860
rect 18334 28806 18336 28858
rect 18398 28806 18410 28858
rect 18472 28806 18474 28858
rect 18312 28804 18336 28806
rect 18392 28804 18416 28806
rect 18472 28804 18496 28806
rect 18256 28784 18552 28804
rect 21256 28860 21552 28880
rect 21312 28858 21336 28860
rect 21392 28858 21416 28860
rect 21472 28858 21496 28860
rect 21334 28806 21336 28858
rect 21398 28806 21410 28858
rect 21472 28806 21474 28858
rect 21312 28804 21336 28806
rect 21392 28804 21416 28806
rect 21472 28804 21496 28806
rect 21256 28784 21552 28804
rect 24256 28860 24552 28880
rect 24312 28858 24336 28860
rect 24392 28858 24416 28860
rect 24472 28858 24496 28860
rect 24334 28806 24336 28858
rect 24398 28806 24410 28858
rect 24472 28806 24474 28858
rect 24312 28804 24336 28806
rect 24392 28804 24416 28806
rect 24472 28804 24496 28806
rect 24256 28784 24552 28804
rect 1756 28316 2052 28336
rect 1812 28314 1836 28316
rect 1892 28314 1916 28316
rect 1972 28314 1996 28316
rect 1834 28262 1836 28314
rect 1898 28262 1910 28314
rect 1972 28262 1974 28314
rect 1812 28260 1836 28262
rect 1892 28260 1916 28262
rect 1972 28260 1996 28262
rect 1756 28240 2052 28260
rect 4756 28316 5052 28336
rect 4812 28314 4836 28316
rect 4892 28314 4916 28316
rect 4972 28314 4996 28316
rect 4834 28262 4836 28314
rect 4898 28262 4910 28314
rect 4972 28262 4974 28314
rect 4812 28260 4836 28262
rect 4892 28260 4916 28262
rect 4972 28260 4996 28262
rect 4756 28240 5052 28260
rect 7756 28316 8052 28336
rect 7812 28314 7836 28316
rect 7892 28314 7916 28316
rect 7972 28314 7996 28316
rect 7834 28262 7836 28314
rect 7898 28262 7910 28314
rect 7972 28262 7974 28314
rect 7812 28260 7836 28262
rect 7892 28260 7916 28262
rect 7972 28260 7996 28262
rect 7756 28240 8052 28260
rect 10756 28316 11052 28336
rect 10812 28314 10836 28316
rect 10892 28314 10916 28316
rect 10972 28314 10996 28316
rect 10834 28262 10836 28314
rect 10898 28262 10910 28314
rect 10972 28262 10974 28314
rect 10812 28260 10836 28262
rect 10892 28260 10916 28262
rect 10972 28260 10996 28262
rect 10756 28240 11052 28260
rect 13756 28316 14052 28336
rect 13812 28314 13836 28316
rect 13892 28314 13916 28316
rect 13972 28314 13996 28316
rect 13834 28262 13836 28314
rect 13898 28262 13910 28314
rect 13972 28262 13974 28314
rect 13812 28260 13836 28262
rect 13892 28260 13916 28262
rect 13972 28260 13996 28262
rect 13756 28240 14052 28260
rect 16756 28316 17052 28336
rect 16812 28314 16836 28316
rect 16892 28314 16916 28316
rect 16972 28314 16996 28316
rect 16834 28262 16836 28314
rect 16898 28262 16910 28314
rect 16972 28262 16974 28314
rect 16812 28260 16836 28262
rect 16892 28260 16916 28262
rect 16972 28260 16996 28262
rect 16756 28240 17052 28260
rect 19756 28316 20052 28336
rect 19812 28314 19836 28316
rect 19892 28314 19916 28316
rect 19972 28314 19996 28316
rect 19834 28262 19836 28314
rect 19898 28262 19910 28314
rect 19972 28262 19974 28314
rect 19812 28260 19836 28262
rect 19892 28260 19916 28262
rect 19972 28260 19996 28262
rect 19756 28240 20052 28260
rect 22756 28316 23052 28336
rect 22812 28314 22836 28316
rect 22892 28314 22916 28316
rect 22972 28314 22996 28316
rect 22834 28262 22836 28314
rect 22898 28262 22910 28314
rect 22972 28262 22974 28314
rect 22812 28260 22836 28262
rect 22892 28260 22916 28262
rect 22972 28260 22996 28262
rect 22756 28240 23052 28260
rect 3256 27772 3552 27792
rect 3312 27770 3336 27772
rect 3392 27770 3416 27772
rect 3472 27770 3496 27772
rect 3334 27718 3336 27770
rect 3398 27718 3410 27770
rect 3472 27718 3474 27770
rect 3312 27716 3336 27718
rect 3392 27716 3416 27718
rect 3472 27716 3496 27718
rect 3256 27696 3552 27716
rect 6256 27772 6552 27792
rect 6312 27770 6336 27772
rect 6392 27770 6416 27772
rect 6472 27770 6496 27772
rect 6334 27718 6336 27770
rect 6398 27718 6410 27770
rect 6472 27718 6474 27770
rect 6312 27716 6336 27718
rect 6392 27716 6416 27718
rect 6472 27716 6496 27718
rect 6256 27696 6552 27716
rect 9256 27772 9552 27792
rect 9312 27770 9336 27772
rect 9392 27770 9416 27772
rect 9472 27770 9496 27772
rect 9334 27718 9336 27770
rect 9398 27718 9410 27770
rect 9472 27718 9474 27770
rect 9312 27716 9336 27718
rect 9392 27716 9416 27718
rect 9472 27716 9496 27718
rect 9256 27696 9552 27716
rect 12256 27772 12552 27792
rect 12312 27770 12336 27772
rect 12392 27770 12416 27772
rect 12472 27770 12496 27772
rect 12334 27718 12336 27770
rect 12398 27718 12410 27770
rect 12472 27718 12474 27770
rect 12312 27716 12336 27718
rect 12392 27716 12416 27718
rect 12472 27716 12496 27718
rect 12256 27696 12552 27716
rect 15256 27772 15552 27792
rect 15312 27770 15336 27772
rect 15392 27770 15416 27772
rect 15472 27770 15496 27772
rect 15334 27718 15336 27770
rect 15398 27718 15410 27770
rect 15472 27718 15474 27770
rect 15312 27716 15336 27718
rect 15392 27716 15416 27718
rect 15472 27716 15496 27718
rect 15256 27696 15552 27716
rect 18256 27772 18552 27792
rect 18312 27770 18336 27772
rect 18392 27770 18416 27772
rect 18472 27770 18496 27772
rect 18334 27718 18336 27770
rect 18398 27718 18410 27770
rect 18472 27718 18474 27770
rect 18312 27716 18336 27718
rect 18392 27716 18416 27718
rect 18472 27716 18496 27718
rect 18256 27696 18552 27716
rect 21256 27772 21552 27792
rect 21312 27770 21336 27772
rect 21392 27770 21416 27772
rect 21472 27770 21496 27772
rect 21334 27718 21336 27770
rect 21398 27718 21410 27770
rect 21472 27718 21474 27770
rect 21312 27716 21336 27718
rect 21392 27716 21416 27718
rect 21472 27716 21496 27718
rect 21256 27696 21552 27716
rect 24256 27772 24552 27792
rect 24312 27770 24336 27772
rect 24392 27770 24416 27772
rect 24472 27770 24496 27772
rect 24334 27718 24336 27770
rect 24398 27718 24410 27770
rect 24472 27718 24474 27770
rect 24312 27716 24336 27718
rect 24392 27716 24416 27718
rect 24472 27716 24496 27718
rect 24256 27696 24552 27716
rect 24596 27470 24624 30926
rect 24858 30871 24914 30926
rect 25756 29404 26052 29424
rect 25812 29402 25836 29404
rect 25892 29402 25916 29404
rect 25972 29402 25996 29404
rect 25834 29350 25836 29402
rect 25898 29350 25910 29402
rect 25972 29350 25974 29402
rect 25812 29348 25836 29350
rect 25892 29348 25916 29350
rect 25972 29348 25996 29350
rect 25756 29328 26052 29348
rect 27256 28860 27552 28880
rect 27312 28858 27336 28860
rect 27392 28858 27416 28860
rect 27472 28858 27496 28860
rect 27334 28806 27336 28858
rect 27398 28806 27410 28858
rect 27472 28806 27474 28858
rect 27312 28804 27336 28806
rect 27392 28804 27416 28806
rect 27472 28804 27496 28806
rect 27256 28784 27552 28804
rect 25756 28316 26052 28336
rect 25812 28314 25836 28316
rect 25892 28314 25916 28316
rect 25972 28314 25996 28316
rect 25834 28262 25836 28314
rect 25898 28262 25910 28314
rect 25972 28262 25974 28314
rect 25812 28260 25836 28262
rect 25892 28260 25916 28262
rect 25972 28260 25996 28262
rect 25756 28240 26052 28260
rect 27256 27772 27552 27792
rect 27312 27770 27336 27772
rect 27392 27770 27416 27772
rect 27472 27770 27496 27772
rect 27334 27718 27336 27770
rect 27398 27718 27410 27770
rect 27472 27718 27474 27770
rect 27312 27716 27336 27718
rect 27392 27716 27416 27718
rect 27472 27716 27496 27718
rect 27256 27696 27552 27716
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 23112 27396 23164 27402
rect 23112 27338 23164 27344
rect 1756 27228 2052 27248
rect 1812 27226 1836 27228
rect 1892 27226 1916 27228
rect 1972 27226 1996 27228
rect 1834 27174 1836 27226
rect 1898 27174 1910 27226
rect 1972 27174 1974 27226
rect 1812 27172 1836 27174
rect 1892 27172 1916 27174
rect 1972 27172 1996 27174
rect 1756 27152 2052 27172
rect 4756 27228 5052 27248
rect 4812 27226 4836 27228
rect 4892 27226 4916 27228
rect 4972 27226 4996 27228
rect 4834 27174 4836 27226
rect 4898 27174 4910 27226
rect 4972 27174 4974 27226
rect 4812 27172 4836 27174
rect 4892 27172 4916 27174
rect 4972 27172 4996 27174
rect 4756 27152 5052 27172
rect 7756 27228 8052 27248
rect 7812 27226 7836 27228
rect 7892 27226 7916 27228
rect 7972 27226 7996 27228
rect 7834 27174 7836 27226
rect 7898 27174 7910 27226
rect 7972 27174 7974 27226
rect 7812 27172 7836 27174
rect 7892 27172 7916 27174
rect 7972 27172 7996 27174
rect 7756 27152 8052 27172
rect 10756 27228 11052 27248
rect 10812 27226 10836 27228
rect 10892 27226 10916 27228
rect 10972 27226 10996 27228
rect 10834 27174 10836 27226
rect 10898 27174 10910 27226
rect 10972 27174 10974 27226
rect 10812 27172 10836 27174
rect 10892 27172 10916 27174
rect 10972 27172 10996 27174
rect 10756 27152 11052 27172
rect 13756 27228 14052 27248
rect 13812 27226 13836 27228
rect 13892 27226 13916 27228
rect 13972 27226 13996 27228
rect 13834 27174 13836 27226
rect 13898 27174 13910 27226
rect 13972 27174 13974 27226
rect 13812 27172 13836 27174
rect 13892 27172 13916 27174
rect 13972 27172 13996 27174
rect 13756 27152 14052 27172
rect 16756 27228 17052 27248
rect 16812 27226 16836 27228
rect 16892 27226 16916 27228
rect 16972 27226 16996 27228
rect 16834 27174 16836 27226
rect 16898 27174 16910 27226
rect 16972 27174 16974 27226
rect 16812 27172 16836 27174
rect 16892 27172 16916 27174
rect 16972 27172 16996 27174
rect 16756 27152 17052 27172
rect 19756 27228 20052 27248
rect 19812 27226 19836 27228
rect 19892 27226 19916 27228
rect 19972 27226 19996 27228
rect 19834 27174 19836 27226
rect 19898 27174 19910 27226
rect 19972 27174 19974 27226
rect 19812 27172 19836 27174
rect 19892 27172 19916 27174
rect 19972 27172 19996 27174
rect 19756 27152 20052 27172
rect 22756 27228 23052 27248
rect 22812 27226 22836 27228
rect 22892 27226 22916 27228
rect 22972 27226 22996 27228
rect 22834 27174 22836 27226
rect 22898 27174 22910 27226
rect 22972 27174 22974 27226
rect 22812 27172 22836 27174
rect 22892 27172 22916 27174
rect 22972 27172 22996 27174
rect 22756 27152 23052 27172
rect 3256 26684 3552 26704
rect 3312 26682 3336 26684
rect 3392 26682 3416 26684
rect 3472 26682 3496 26684
rect 3334 26630 3336 26682
rect 3398 26630 3410 26682
rect 3472 26630 3474 26682
rect 3312 26628 3336 26630
rect 3392 26628 3416 26630
rect 3472 26628 3496 26630
rect 3256 26608 3552 26628
rect 6256 26684 6552 26704
rect 6312 26682 6336 26684
rect 6392 26682 6416 26684
rect 6472 26682 6496 26684
rect 6334 26630 6336 26682
rect 6398 26630 6410 26682
rect 6472 26630 6474 26682
rect 6312 26628 6336 26630
rect 6392 26628 6416 26630
rect 6472 26628 6496 26630
rect 6256 26608 6552 26628
rect 9256 26684 9552 26704
rect 9312 26682 9336 26684
rect 9392 26682 9416 26684
rect 9472 26682 9496 26684
rect 9334 26630 9336 26682
rect 9398 26630 9410 26682
rect 9472 26630 9474 26682
rect 9312 26628 9336 26630
rect 9392 26628 9416 26630
rect 9472 26628 9496 26630
rect 9256 26608 9552 26628
rect 12256 26684 12552 26704
rect 12312 26682 12336 26684
rect 12392 26682 12416 26684
rect 12472 26682 12496 26684
rect 12334 26630 12336 26682
rect 12398 26630 12410 26682
rect 12472 26630 12474 26682
rect 12312 26628 12336 26630
rect 12392 26628 12416 26630
rect 12472 26628 12496 26630
rect 12256 26608 12552 26628
rect 15256 26684 15552 26704
rect 15312 26682 15336 26684
rect 15392 26682 15416 26684
rect 15472 26682 15496 26684
rect 15334 26630 15336 26682
rect 15398 26630 15410 26682
rect 15472 26630 15474 26682
rect 15312 26628 15336 26630
rect 15392 26628 15416 26630
rect 15472 26628 15496 26630
rect 15256 26608 15552 26628
rect 18256 26684 18552 26704
rect 18312 26682 18336 26684
rect 18392 26682 18416 26684
rect 18472 26682 18496 26684
rect 18334 26630 18336 26682
rect 18398 26630 18410 26682
rect 18472 26630 18474 26682
rect 18312 26628 18336 26630
rect 18392 26628 18416 26630
rect 18472 26628 18496 26630
rect 18256 26608 18552 26628
rect 21256 26684 21552 26704
rect 21312 26682 21336 26684
rect 21392 26682 21416 26684
rect 21472 26682 21496 26684
rect 21334 26630 21336 26682
rect 21398 26630 21410 26682
rect 21472 26630 21474 26682
rect 21312 26628 21336 26630
rect 21392 26628 21416 26630
rect 21472 26628 21496 26630
rect 21256 26608 21552 26628
rect 1756 26140 2052 26160
rect 1812 26138 1836 26140
rect 1892 26138 1916 26140
rect 1972 26138 1996 26140
rect 1834 26086 1836 26138
rect 1898 26086 1910 26138
rect 1972 26086 1974 26138
rect 1812 26084 1836 26086
rect 1892 26084 1916 26086
rect 1972 26084 1996 26086
rect 1756 26064 2052 26084
rect 4756 26140 5052 26160
rect 4812 26138 4836 26140
rect 4892 26138 4916 26140
rect 4972 26138 4996 26140
rect 4834 26086 4836 26138
rect 4898 26086 4910 26138
rect 4972 26086 4974 26138
rect 4812 26084 4836 26086
rect 4892 26084 4916 26086
rect 4972 26084 4996 26086
rect 4756 26064 5052 26084
rect 7756 26140 8052 26160
rect 7812 26138 7836 26140
rect 7892 26138 7916 26140
rect 7972 26138 7996 26140
rect 7834 26086 7836 26138
rect 7898 26086 7910 26138
rect 7972 26086 7974 26138
rect 7812 26084 7836 26086
rect 7892 26084 7916 26086
rect 7972 26084 7996 26086
rect 7756 26064 8052 26084
rect 10756 26140 11052 26160
rect 10812 26138 10836 26140
rect 10892 26138 10916 26140
rect 10972 26138 10996 26140
rect 10834 26086 10836 26138
rect 10898 26086 10910 26138
rect 10972 26086 10974 26138
rect 10812 26084 10836 26086
rect 10892 26084 10916 26086
rect 10972 26084 10996 26086
rect 10756 26064 11052 26084
rect 13756 26140 14052 26160
rect 13812 26138 13836 26140
rect 13892 26138 13916 26140
rect 13972 26138 13996 26140
rect 13834 26086 13836 26138
rect 13898 26086 13910 26138
rect 13972 26086 13974 26138
rect 13812 26084 13836 26086
rect 13892 26084 13916 26086
rect 13972 26084 13996 26086
rect 13756 26064 14052 26084
rect 16756 26140 17052 26160
rect 16812 26138 16836 26140
rect 16892 26138 16916 26140
rect 16972 26138 16996 26140
rect 16834 26086 16836 26138
rect 16898 26086 16910 26138
rect 16972 26086 16974 26138
rect 16812 26084 16836 26086
rect 16892 26084 16916 26086
rect 16972 26084 16996 26086
rect 16756 26064 17052 26084
rect 19756 26140 20052 26160
rect 19812 26138 19836 26140
rect 19892 26138 19916 26140
rect 19972 26138 19996 26140
rect 19834 26086 19836 26138
rect 19898 26086 19910 26138
rect 19972 26086 19974 26138
rect 19812 26084 19836 26086
rect 19892 26084 19916 26086
rect 19972 26084 19996 26086
rect 19756 26064 20052 26084
rect 22756 26140 23052 26160
rect 22812 26138 22836 26140
rect 22892 26138 22916 26140
rect 22972 26138 22996 26140
rect 22834 26086 22836 26138
rect 22898 26086 22910 26138
rect 22972 26086 22974 26138
rect 22812 26084 22836 26086
rect 22892 26084 22916 26086
rect 22972 26084 22996 26086
rect 22756 26064 23052 26084
rect 3256 25596 3552 25616
rect 3312 25594 3336 25596
rect 3392 25594 3416 25596
rect 3472 25594 3496 25596
rect 3334 25542 3336 25594
rect 3398 25542 3410 25594
rect 3472 25542 3474 25594
rect 3312 25540 3336 25542
rect 3392 25540 3416 25542
rect 3472 25540 3496 25542
rect 3256 25520 3552 25540
rect 6256 25596 6552 25616
rect 6312 25594 6336 25596
rect 6392 25594 6416 25596
rect 6472 25594 6496 25596
rect 6334 25542 6336 25594
rect 6398 25542 6410 25594
rect 6472 25542 6474 25594
rect 6312 25540 6336 25542
rect 6392 25540 6416 25542
rect 6472 25540 6496 25542
rect 6256 25520 6552 25540
rect 9256 25596 9552 25616
rect 9312 25594 9336 25596
rect 9392 25594 9416 25596
rect 9472 25594 9496 25596
rect 9334 25542 9336 25594
rect 9398 25542 9410 25594
rect 9472 25542 9474 25594
rect 9312 25540 9336 25542
rect 9392 25540 9416 25542
rect 9472 25540 9496 25542
rect 9256 25520 9552 25540
rect 12256 25596 12552 25616
rect 12312 25594 12336 25596
rect 12392 25594 12416 25596
rect 12472 25594 12496 25596
rect 12334 25542 12336 25594
rect 12398 25542 12410 25594
rect 12472 25542 12474 25594
rect 12312 25540 12336 25542
rect 12392 25540 12416 25542
rect 12472 25540 12496 25542
rect 12256 25520 12552 25540
rect 15256 25596 15552 25616
rect 15312 25594 15336 25596
rect 15392 25594 15416 25596
rect 15472 25594 15496 25596
rect 15334 25542 15336 25594
rect 15398 25542 15410 25594
rect 15472 25542 15474 25594
rect 15312 25540 15336 25542
rect 15392 25540 15416 25542
rect 15472 25540 15496 25542
rect 15256 25520 15552 25540
rect 18256 25596 18552 25616
rect 18312 25594 18336 25596
rect 18392 25594 18416 25596
rect 18472 25594 18496 25596
rect 18334 25542 18336 25594
rect 18398 25542 18410 25594
rect 18472 25542 18474 25594
rect 18312 25540 18336 25542
rect 18392 25540 18416 25542
rect 18472 25540 18496 25542
rect 18256 25520 18552 25540
rect 21256 25596 21552 25616
rect 21312 25594 21336 25596
rect 21392 25594 21416 25596
rect 21472 25594 21496 25596
rect 21334 25542 21336 25594
rect 21398 25542 21410 25594
rect 21472 25542 21474 25594
rect 21312 25540 21336 25542
rect 21392 25540 21416 25542
rect 21472 25540 21496 25542
rect 21256 25520 21552 25540
rect 1756 25052 2052 25072
rect 1812 25050 1836 25052
rect 1892 25050 1916 25052
rect 1972 25050 1996 25052
rect 1834 24998 1836 25050
rect 1898 24998 1910 25050
rect 1972 24998 1974 25050
rect 1812 24996 1836 24998
rect 1892 24996 1916 24998
rect 1972 24996 1996 24998
rect 1756 24976 2052 24996
rect 4756 25052 5052 25072
rect 4812 25050 4836 25052
rect 4892 25050 4916 25052
rect 4972 25050 4996 25052
rect 4834 24998 4836 25050
rect 4898 24998 4910 25050
rect 4972 24998 4974 25050
rect 4812 24996 4836 24998
rect 4892 24996 4916 24998
rect 4972 24996 4996 24998
rect 4756 24976 5052 24996
rect 7756 25052 8052 25072
rect 7812 25050 7836 25052
rect 7892 25050 7916 25052
rect 7972 25050 7996 25052
rect 7834 24998 7836 25050
rect 7898 24998 7910 25050
rect 7972 24998 7974 25050
rect 7812 24996 7836 24998
rect 7892 24996 7916 24998
rect 7972 24996 7996 24998
rect 7756 24976 8052 24996
rect 10756 25052 11052 25072
rect 10812 25050 10836 25052
rect 10892 25050 10916 25052
rect 10972 25050 10996 25052
rect 10834 24998 10836 25050
rect 10898 24998 10910 25050
rect 10972 24998 10974 25050
rect 10812 24996 10836 24998
rect 10892 24996 10916 24998
rect 10972 24996 10996 24998
rect 10756 24976 11052 24996
rect 13756 25052 14052 25072
rect 13812 25050 13836 25052
rect 13892 25050 13916 25052
rect 13972 25050 13996 25052
rect 13834 24998 13836 25050
rect 13898 24998 13910 25050
rect 13972 24998 13974 25050
rect 13812 24996 13836 24998
rect 13892 24996 13916 24998
rect 13972 24996 13996 24998
rect 13756 24976 14052 24996
rect 16756 25052 17052 25072
rect 16812 25050 16836 25052
rect 16892 25050 16916 25052
rect 16972 25050 16996 25052
rect 16834 24998 16836 25050
rect 16898 24998 16910 25050
rect 16972 24998 16974 25050
rect 16812 24996 16836 24998
rect 16892 24996 16916 24998
rect 16972 24996 16996 24998
rect 16756 24976 17052 24996
rect 19756 25052 20052 25072
rect 19812 25050 19836 25052
rect 19892 25050 19916 25052
rect 19972 25050 19996 25052
rect 19834 24998 19836 25050
rect 19898 24998 19910 25050
rect 19972 24998 19974 25050
rect 19812 24996 19836 24998
rect 19892 24996 19916 24998
rect 19972 24996 19996 24998
rect 19756 24976 20052 24996
rect 22756 25052 23052 25072
rect 22812 25050 22836 25052
rect 22892 25050 22916 25052
rect 22972 25050 22996 25052
rect 22834 24998 22836 25050
rect 22898 24998 22910 25050
rect 22972 24998 22974 25050
rect 22812 24996 22836 24998
rect 22892 24996 22916 24998
rect 22972 24996 22996 24998
rect 22756 24976 23052 24996
rect 3256 24508 3552 24528
rect 3312 24506 3336 24508
rect 3392 24506 3416 24508
rect 3472 24506 3496 24508
rect 3334 24454 3336 24506
rect 3398 24454 3410 24506
rect 3472 24454 3474 24506
rect 3312 24452 3336 24454
rect 3392 24452 3416 24454
rect 3472 24452 3496 24454
rect 3256 24432 3552 24452
rect 6256 24508 6552 24528
rect 6312 24506 6336 24508
rect 6392 24506 6416 24508
rect 6472 24506 6496 24508
rect 6334 24454 6336 24506
rect 6398 24454 6410 24506
rect 6472 24454 6474 24506
rect 6312 24452 6336 24454
rect 6392 24452 6416 24454
rect 6472 24452 6496 24454
rect 6256 24432 6552 24452
rect 9256 24508 9552 24528
rect 9312 24506 9336 24508
rect 9392 24506 9416 24508
rect 9472 24506 9496 24508
rect 9334 24454 9336 24506
rect 9398 24454 9410 24506
rect 9472 24454 9474 24506
rect 9312 24452 9336 24454
rect 9392 24452 9416 24454
rect 9472 24452 9496 24454
rect 9256 24432 9552 24452
rect 12256 24508 12552 24528
rect 12312 24506 12336 24508
rect 12392 24506 12416 24508
rect 12472 24506 12496 24508
rect 12334 24454 12336 24506
rect 12398 24454 12410 24506
rect 12472 24454 12474 24506
rect 12312 24452 12336 24454
rect 12392 24452 12416 24454
rect 12472 24452 12496 24454
rect 12256 24432 12552 24452
rect 15256 24508 15552 24528
rect 15312 24506 15336 24508
rect 15392 24506 15416 24508
rect 15472 24506 15496 24508
rect 15334 24454 15336 24506
rect 15398 24454 15410 24506
rect 15472 24454 15474 24506
rect 15312 24452 15336 24454
rect 15392 24452 15416 24454
rect 15472 24452 15496 24454
rect 15256 24432 15552 24452
rect 18256 24508 18552 24528
rect 18312 24506 18336 24508
rect 18392 24506 18416 24508
rect 18472 24506 18496 24508
rect 18334 24454 18336 24506
rect 18398 24454 18410 24506
rect 18472 24454 18474 24506
rect 18312 24452 18336 24454
rect 18392 24452 18416 24454
rect 18472 24452 18496 24454
rect 18256 24432 18552 24452
rect 21256 24508 21552 24528
rect 21312 24506 21336 24508
rect 21392 24506 21416 24508
rect 21472 24506 21496 24508
rect 21334 24454 21336 24506
rect 21398 24454 21410 24506
rect 21472 24454 21474 24506
rect 21312 24452 21336 24454
rect 21392 24452 21416 24454
rect 21472 24452 21496 24454
rect 21256 24432 21552 24452
rect 1756 23964 2052 23984
rect 1812 23962 1836 23964
rect 1892 23962 1916 23964
rect 1972 23962 1996 23964
rect 1834 23910 1836 23962
rect 1898 23910 1910 23962
rect 1972 23910 1974 23962
rect 1812 23908 1836 23910
rect 1892 23908 1916 23910
rect 1972 23908 1996 23910
rect 1756 23888 2052 23908
rect 4756 23964 5052 23984
rect 4812 23962 4836 23964
rect 4892 23962 4916 23964
rect 4972 23962 4996 23964
rect 4834 23910 4836 23962
rect 4898 23910 4910 23962
rect 4972 23910 4974 23962
rect 4812 23908 4836 23910
rect 4892 23908 4916 23910
rect 4972 23908 4996 23910
rect 4756 23888 5052 23908
rect 7756 23964 8052 23984
rect 7812 23962 7836 23964
rect 7892 23962 7916 23964
rect 7972 23962 7996 23964
rect 7834 23910 7836 23962
rect 7898 23910 7910 23962
rect 7972 23910 7974 23962
rect 7812 23908 7836 23910
rect 7892 23908 7916 23910
rect 7972 23908 7996 23910
rect 7756 23888 8052 23908
rect 10756 23964 11052 23984
rect 10812 23962 10836 23964
rect 10892 23962 10916 23964
rect 10972 23962 10996 23964
rect 10834 23910 10836 23962
rect 10898 23910 10910 23962
rect 10972 23910 10974 23962
rect 10812 23908 10836 23910
rect 10892 23908 10916 23910
rect 10972 23908 10996 23910
rect 10756 23888 11052 23908
rect 13756 23964 14052 23984
rect 13812 23962 13836 23964
rect 13892 23962 13916 23964
rect 13972 23962 13996 23964
rect 13834 23910 13836 23962
rect 13898 23910 13910 23962
rect 13972 23910 13974 23962
rect 13812 23908 13836 23910
rect 13892 23908 13916 23910
rect 13972 23908 13996 23910
rect 13756 23888 14052 23908
rect 16756 23964 17052 23984
rect 16812 23962 16836 23964
rect 16892 23962 16916 23964
rect 16972 23962 16996 23964
rect 16834 23910 16836 23962
rect 16898 23910 16910 23962
rect 16972 23910 16974 23962
rect 16812 23908 16836 23910
rect 16892 23908 16916 23910
rect 16972 23908 16996 23910
rect 16756 23888 17052 23908
rect 19756 23964 20052 23984
rect 19812 23962 19836 23964
rect 19892 23962 19916 23964
rect 19972 23962 19996 23964
rect 19834 23910 19836 23962
rect 19898 23910 19910 23962
rect 19972 23910 19974 23962
rect 19812 23908 19836 23910
rect 19892 23908 19916 23910
rect 19972 23908 19996 23910
rect 19756 23888 20052 23908
rect 22756 23964 23052 23984
rect 22812 23962 22836 23964
rect 22892 23962 22916 23964
rect 22972 23962 22996 23964
rect 22834 23910 22836 23962
rect 22898 23910 22910 23962
rect 22972 23910 22974 23962
rect 22812 23908 22836 23910
rect 22892 23908 22916 23910
rect 22972 23908 22996 23910
rect 22756 23888 23052 23908
rect 3256 23420 3552 23440
rect 3312 23418 3336 23420
rect 3392 23418 3416 23420
rect 3472 23418 3496 23420
rect 3334 23366 3336 23418
rect 3398 23366 3410 23418
rect 3472 23366 3474 23418
rect 3312 23364 3336 23366
rect 3392 23364 3416 23366
rect 3472 23364 3496 23366
rect 3256 23344 3552 23364
rect 6256 23420 6552 23440
rect 6312 23418 6336 23420
rect 6392 23418 6416 23420
rect 6472 23418 6496 23420
rect 6334 23366 6336 23418
rect 6398 23366 6410 23418
rect 6472 23366 6474 23418
rect 6312 23364 6336 23366
rect 6392 23364 6416 23366
rect 6472 23364 6496 23366
rect 6256 23344 6552 23364
rect 9256 23420 9552 23440
rect 9312 23418 9336 23420
rect 9392 23418 9416 23420
rect 9472 23418 9496 23420
rect 9334 23366 9336 23418
rect 9398 23366 9410 23418
rect 9472 23366 9474 23418
rect 9312 23364 9336 23366
rect 9392 23364 9416 23366
rect 9472 23364 9496 23366
rect 9256 23344 9552 23364
rect 12256 23420 12552 23440
rect 12312 23418 12336 23420
rect 12392 23418 12416 23420
rect 12472 23418 12496 23420
rect 12334 23366 12336 23418
rect 12398 23366 12410 23418
rect 12472 23366 12474 23418
rect 12312 23364 12336 23366
rect 12392 23364 12416 23366
rect 12472 23364 12496 23366
rect 12256 23344 12552 23364
rect 15256 23420 15552 23440
rect 15312 23418 15336 23420
rect 15392 23418 15416 23420
rect 15472 23418 15496 23420
rect 15334 23366 15336 23418
rect 15398 23366 15410 23418
rect 15472 23366 15474 23418
rect 15312 23364 15336 23366
rect 15392 23364 15416 23366
rect 15472 23364 15496 23366
rect 15256 23344 15552 23364
rect 18256 23420 18552 23440
rect 18312 23418 18336 23420
rect 18392 23418 18416 23420
rect 18472 23418 18496 23420
rect 18334 23366 18336 23418
rect 18398 23366 18410 23418
rect 18472 23366 18474 23418
rect 18312 23364 18336 23366
rect 18392 23364 18416 23366
rect 18472 23364 18496 23366
rect 18256 23344 18552 23364
rect 21256 23420 21552 23440
rect 21312 23418 21336 23420
rect 21392 23418 21416 23420
rect 21472 23418 21496 23420
rect 21334 23366 21336 23418
rect 21398 23366 21410 23418
rect 21472 23366 21474 23418
rect 21312 23364 21336 23366
rect 21392 23364 21416 23366
rect 21472 23364 21496 23366
rect 21256 23344 21552 23364
rect 1756 22876 2052 22896
rect 1812 22874 1836 22876
rect 1892 22874 1916 22876
rect 1972 22874 1996 22876
rect 1834 22822 1836 22874
rect 1898 22822 1910 22874
rect 1972 22822 1974 22874
rect 1812 22820 1836 22822
rect 1892 22820 1916 22822
rect 1972 22820 1996 22822
rect 1756 22800 2052 22820
rect 4756 22876 5052 22896
rect 4812 22874 4836 22876
rect 4892 22874 4916 22876
rect 4972 22874 4996 22876
rect 4834 22822 4836 22874
rect 4898 22822 4910 22874
rect 4972 22822 4974 22874
rect 4812 22820 4836 22822
rect 4892 22820 4916 22822
rect 4972 22820 4996 22822
rect 4756 22800 5052 22820
rect 7756 22876 8052 22896
rect 7812 22874 7836 22876
rect 7892 22874 7916 22876
rect 7972 22874 7996 22876
rect 7834 22822 7836 22874
rect 7898 22822 7910 22874
rect 7972 22822 7974 22874
rect 7812 22820 7836 22822
rect 7892 22820 7916 22822
rect 7972 22820 7996 22822
rect 7756 22800 8052 22820
rect 10756 22876 11052 22896
rect 10812 22874 10836 22876
rect 10892 22874 10916 22876
rect 10972 22874 10996 22876
rect 10834 22822 10836 22874
rect 10898 22822 10910 22874
rect 10972 22822 10974 22874
rect 10812 22820 10836 22822
rect 10892 22820 10916 22822
rect 10972 22820 10996 22822
rect 10756 22800 11052 22820
rect 13756 22876 14052 22896
rect 13812 22874 13836 22876
rect 13892 22874 13916 22876
rect 13972 22874 13996 22876
rect 13834 22822 13836 22874
rect 13898 22822 13910 22874
rect 13972 22822 13974 22874
rect 13812 22820 13836 22822
rect 13892 22820 13916 22822
rect 13972 22820 13996 22822
rect 13756 22800 14052 22820
rect 16756 22876 17052 22896
rect 16812 22874 16836 22876
rect 16892 22874 16916 22876
rect 16972 22874 16996 22876
rect 16834 22822 16836 22874
rect 16898 22822 16910 22874
rect 16972 22822 16974 22874
rect 16812 22820 16836 22822
rect 16892 22820 16916 22822
rect 16972 22820 16996 22822
rect 16756 22800 17052 22820
rect 19756 22876 20052 22896
rect 19812 22874 19836 22876
rect 19892 22874 19916 22876
rect 19972 22874 19996 22876
rect 19834 22822 19836 22874
rect 19898 22822 19910 22874
rect 19972 22822 19974 22874
rect 19812 22820 19836 22822
rect 19892 22820 19916 22822
rect 19972 22820 19996 22822
rect 19756 22800 20052 22820
rect 22756 22876 23052 22896
rect 22812 22874 22836 22876
rect 22892 22874 22916 22876
rect 22972 22874 22996 22876
rect 22834 22822 22836 22874
rect 22898 22822 22910 22874
rect 22972 22822 22974 22874
rect 22812 22820 22836 22822
rect 22892 22820 22916 22822
rect 22972 22820 22996 22822
rect 22756 22800 23052 22820
rect 3256 22332 3552 22352
rect 3312 22330 3336 22332
rect 3392 22330 3416 22332
rect 3472 22330 3496 22332
rect 3334 22278 3336 22330
rect 3398 22278 3410 22330
rect 3472 22278 3474 22330
rect 3312 22276 3336 22278
rect 3392 22276 3416 22278
rect 3472 22276 3496 22278
rect 3256 22256 3552 22276
rect 6256 22332 6552 22352
rect 6312 22330 6336 22332
rect 6392 22330 6416 22332
rect 6472 22330 6496 22332
rect 6334 22278 6336 22330
rect 6398 22278 6410 22330
rect 6472 22278 6474 22330
rect 6312 22276 6336 22278
rect 6392 22276 6416 22278
rect 6472 22276 6496 22278
rect 6256 22256 6552 22276
rect 9256 22332 9552 22352
rect 9312 22330 9336 22332
rect 9392 22330 9416 22332
rect 9472 22330 9496 22332
rect 9334 22278 9336 22330
rect 9398 22278 9410 22330
rect 9472 22278 9474 22330
rect 9312 22276 9336 22278
rect 9392 22276 9416 22278
rect 9472 22276 9496 22278
rect 9256 22256 9552 22276
rect 12256 22332 12552 22352
rect 12312 22330 12336 22332
rect 12392 22330 12416 22332
rect 12472 22330 12496 22332
rect 12334 22278 12336 22330
rect 12398 22278 12410 22330
rect 12472 22278 12474 22330
rect 12312 22276 12336 22278
rect 12392 22276 12416 22278
rect 12472 22276 12496 22278
rect 12256 22256 12552 22276
rect 15256 22332 15552 22352
rect 15312 22330 15336 22332
rect 15392 22330 15416 22332
rect 15472 22330 15496 22332
rect 15334 22278 15336 22330
rect 15398 22278 15410 22330
rect 15472 22278 15474 22330
rect 15312 22276 15336 22278
rect 15392 22276 15416 22278
rect 15472 22276 15496 22278
rect 15256 22256 15552 22276
rect 18256 22332 18552 22352
rect 18312 22330 18336 22332
rect 18392 22330 18416 22332
rect 18472 22330 18496 22332
rect 18334 22278 18336 22330
rect 18398 22278 18410 22330
rect 18472 22278 18474 22330
rect 18312 22276 18336 22278
rect 18392 22276 18416 22278
rect 18472 22276 18496 22278
rect 18256 22256 18552 22276
rect 21256 22332 21552 22352
rect 21312 22330 21336 22332
rect 21392 22330 21416 22332
rect 21472 22330 21496 22332
rect 21334 22278 21336 22330
rect 21398 22278 21410 22330
rect 21472 22278 21474 22330
rect 21312 22276 21336 22278
rect 21392 22276 21416 22278
rect 21472 22276 21496 22278
rect 21256 22256 21552 22276
rect 1756 21788 2052 21808
rect 1812 21786 1836 21788
rect 1892 21786 1916 21788
rect 1972 21786 1996 21788
rect 1834 21734 1836 21786
rect 1898 21734 1910 21786
rect 1972 21734 1974 21786
rect 1812 21732 1836 21734
rect 1892 21732 1916 21734
rect 1972 21732 1996 21734
rect 1756 21712 2052 21732
rect 4756 21788 5052 21808
rect 4812 21786 4836 21788
rect 4892 21786 4916 21788
rect 4972 21786 4996 21788
rect 4834 21734 4836 21786
rect 4898 21734 4910 21786
rect 4972 21734 4974 21786
rect 4812 21732 4836 21734
rect 4892 21732 4916 21734
rect 4972 21732 4996 21734
rect 4756 21712 5052 21732
rect 7756 21788 8052 21808
rect 7812 21786 7836 21788
rect 7892 21786 7916 21788
rect 7972 21786 7996 21788
rect 7834 21734 7836 21786
rect 7898 21734 7910 21786
rect 7972 21734 7974 21786
rect 7812 21732 7836 21734
rect 7892 21732 7916 21734
rect 7972 21732 7996 21734
rect 7756 21712 8052 21732
rect 10756 21788 11052 21808
rect 10812 21786 10836 21788
rect 10892 21786 10916 21788
rect 10972 21786 10996 21788
rect 10834 21734 10836 21786
rect 10898 21734 10910 21786
rect 10972 21734 10974 21786
rect 10812 21732 10836 21734
rect 10892 21732 10916 21734
rect 10972 21732 10996 21734
rect 10756 21712 11052 21732
rect 13756 21788 14052 21808
rect 13812 21786 13836 21788
rect 13892 21786 13916 21788
rect 13972 21786 13996 21788
rect 13834 21734 13836 21786
rect 13898 21734 13910 21786
rect 13972 21734 13974 21786
rect 13812 21732 13836 21734
rect 13892 21732 13916 21734
rect 13972 21732 13996 21734
rect 13756 21712 14052 21732
rect 16756 21788 17052 21808
rect 16812 21786 16836 21788
rect 16892 21786 16916 21788
rect 16972 21786 16996 21788
rect 16834 21734 16836 21786
rect 16898 21734 16910 21786
rect 16972 21734 16974 21786
rect 16812 21732 16836 21734
rect 16892 21732 16916 21734
rect 16972 21732 16996 21734
rect 16756 21712 17052 21732
rect 19756 21788 20052 21808
rect 19812 21786 19836 21788
rect 19892 21786 19916 21788
rect 19972 21786 19996 21788
rect 19834 21734 19836 21786
rect 19898 21734 19910 21786
rect 19972 21734 19974 21786
rect 19812 21732 19836 21734
rect 19892 21732 19916 21734
rect 19972 21732 19996 21734
rect 19756 21712 20052 21732
rect 22756 21788 23052 21808
rect 22812 21786 22836 21788
rect 22892 21786 22916 21788
rect 22972 21786 22996 21788
rect 22834 21734 22836 21786
rect 22898 21734 22910 21786
rect 22972 21734 22974 21786
rect 22812 21732 22836 21734
rect 22892 21732 22916 21734
rect 22972 21732 22996 21734
rect 22756 21712 23052 21732
rect 3256 21244 3552 21264
rect 3312 21242 3336 21244
rect 3392 21242 3416 21244
rect 3472 21242 3496 21244
rect 3334 21190 3336 21242
rect 3398 21190 3410 21242
rect 3472 21190 3474 21242
rect 3312 21188 3336 21190
rect 3392 21188 3416 21190
rect 3472 21188 3496 21190
rect 3256 21168 3552 21188
rect 6256 21244 6552 21264
rect 6312 21242 6336 21244
rect 6392 21242 6416 21244
rect 6472 21242 6496 21244
rect 6334 21190 6336 21242
rect 6398 21190 6410 21242
rect 6472 21190 6474 21242
rect 6312 21188 6336 21190
rect 6392 21188 6416 21190
rect 6472 21188 6496 21190
rect 6256 21168 6552 21188
rect 9256 21244 9552 21264
rect 9312 21242 9336 21244
rect 9392 21242 9416 21244
rect 9472 21242 9496 21244
rect 9334 21190 9336 21242
rect 9398 21190 9410 21242
rect 9472 21190 9474 21242
rect 9312 21188 9336 21190
rect 9392 21188 9416 21190
rect 9472 21188 9496 21190
rect 9256 21168 9552 21188
rect 12256 21244 12552 21264
rect 12312 21242 12336 21244
rect 12392 21242 12416 21244
rect 12472 21242 12496 21244
rect 12334 21190 12336 21242
rect 12398 21190 12410 21242
rect 12472 21190 12474 21242
rect 12312 21188 12336 21190
rect 12392 21188 12416 21190
rect 12472 21188 12496 21190
rect 12256 21168 12552 21188
rect 15256 21244 15552 21264
rect 15312 21242 15336 21244
rect 15392 21242 15416 21244
rect 15472 21242 15496 21244
rect 15334 21190 15336 21242
rect 15398 21190 15410 21242
rect 15472 21190 15474 21242
rect 15312 21188 15336 21190
rect 15392 21188 15416 21190
rect 15472 21188 15496 21190
rect 15256 21168 15552 21188
rect 18256 21244 18552 21264
rect 18312 21242 18336 21244
rect 18392 21242 18416 21244
rect 18472 21242 18496 21244
rect 18334 21190 18336 21242
rect 18398 21190 18410 21242
rect 18472 21190 18474 21242
rect 18312 21188 18336 21190
rect 18392 21188 18416 21190
rect 18472 21188 18496 21190
rect 18256 21168 18552 21188
rect 21256 21244 21552 21264
rect 21312 21242 21336 21244
rect 21392 21242 21416 21244
rect 21472 21242 21496 21244
rect 21334 21190 21336 21242
rect 21398 21190 21410 21242
rect 21472 21190 21474 21242
rect 21312 21188 21336 21190
rect 21392 21188 21416 21190
rect 21472 21188 21496 21190
rect 21256 21168 21552 21188
rect 1756 20700 2052 20720
rect 1812 20698 1836 20700
rect 1892 20698 1916 20700
rect 1972 20698 1996 20700
rect 1834 20646 1836 20698
rect 1898 20646 1910 20698
rect 1972 20646 1974 20698
rect 1812 20644 1836 20646
rect 1892 20644 1916 20646
rect 1972 20644 1996 20646
rect 1756 20624 2052 20644
rect 4756 20700 5052 20720
rect 4812 20698 4836 20700
rect 4892 20698 4916 20700
rect 4972 20698 4996 20700
rect 4834 20646 4836 20698
rect 4898 20646 4910 20698
rect 4972 20646 4974 20698
rect 4812 20644 4836 20646
rect 4892 20644 4916 20646
rect 4972 20644 4996 20646
rect 4756 20624 5052 20644
rect 7756 20700 8052 20720
rect 7812 20698 7836 20700
rect 7892 20698 7916 20700
rect 7972 20698 7996 20700
rect 7834 20646 7836 20698
rect 7898 20646 7910 20698
rect 7972 20646 7974 20698
rect 7812 20644 7836 20646
rect 7892 20644 7916 20646
rect 7972 20644 7996 20646
rect 7756 20624 8052 20644
rect 10756 20700 11052 20720
rect 10812 20698 10836 20700
rect 10892 20698 10916 20700
rect 10972 20698 10996 20700
rect 10834 20646 10836 20698
rect 10898 20646 10910 20698
rect 10972 20646 10974 20698
rect 10812 20644 10836 20646
rect 10892 20644 10916 20646
rect 10972 20644 10996 20646
rect 10756 20624 11052 20644
rect 13756 20700 14052 20720
rect 13812 20698 13836 20700
rect 13892 20698 13916 20700
rect 13972 20698 13996 20700
rect 13834 20646 13836 20698
rect 13898 20646 13910 20698
rect 13972 20646 13974 20698
rect 13812 20644 13836 20646
rect 13892 20644 13916 20646
rect 13972 20644 13996 20646
rect 13756 20624 14052 20644
rect 16756 20700 17052 20720
rect 16812 20698 16836 20700
rect 16892 20698 16916 20700
rect 16972 20698 16996 20700
rect 16834 20646 16836 20698
rect 16898 20646 16910 20698
rect 16972 20646 16974 20698
rect 16812 20644 16836 20646
rect 16892 20644 16916 20646
rect 16972 20644 16996 20646
rect 16756 20624 17052 20644
rect 19756 20700 20052 20720
rect 19812 20698 19836 20700
rect 19892 20698 19916 20700
rect 19972 20698 19996 20700
rect 19834 20646 19836 20698
rect 19898 20646 19910 20698
rect 19972 20646 19974 20698
rect 19812 20644 19836 20646
rect 19892 20644 19916 20646
rect 19972 20644 19996 20646
rect 19756 20624 20052 20644
rect 22756 20700 23052 20720
rect 22812 20698 22836 20700
rect 22892 20698 22916 20700
rect 22972 20698 22996 20700
rect 22834 20646 22836 20698
rect 22898 20646 22910 20698
rect 22972 20646 22974 20698
rect 22812 20644 22836 20646
rect 22892 20644 22916 20646
rect 22972 20644 22996 20646
rect 22756 20624 23052 20644
rect 3256 20156 3552 20176
rect 3312 20154 3336 20156
rect 3392 20154 3416 20156
rect 3472 20154 3496 20156
rect 3334 20102 3336 20154
rect 3398 20102 3410 20154
rect 3472 20102 3474 20154
rect 3312 20100 3336 20102
rect 3392 20100 3416 20102
rect 3472 20100 3496 20102
rect 3256 20080 3552 20100
rect 6256 20156 6552 20176
rect 6312 20154 6336 20156
rect 6392 20154 6416 20156
rect 6472 20154 6496 20156
rect 6334 20102 6336 20154
rect 6398 20102 6410 20154
rect 6472 20102 6474 20154
rect 6312 20100 6336 20102
rect 6392 20100 6416 20102
rect 6472 20100 6496 20102
rect 6256 20080 6552 20100
rect 9256 20156 9552 20176
rect 9312 20154 9336 20156
rect 9392 20154 9416 20156
rect 9472 20154 9496 20156
rect 9334 20102 9336 20154
rect 9398 20102 9410 20154
rect 9472 20102 9474 20154
rect 9312 20100 9336 20102
rect 9392 20100 9416 20102
rect 9472 20100 9496 20102
rect 9256 20080 9552 20100
rect 12256 20156 12552 20176
rect 12312 20154 12336 20156
rect 12392 20154 12416 20156
rect 12472 20154 12496 20156
rect 12334 20102 12336 20154
rect 12398 20102 12410 20154
rect 12472 20102 12474 20154
rect 12312 20100 12336 20102
rect 12392 20100 12416 20102
rect 12472 20100 12496 20102
rect 12256 20080 12552 20100
rect 15256 20156 15552 20176
rect 15312 20154 15336 20156
rect 15392 20154 15416 20156
rect 15472 20154 15496 20156
rect 15334 20102 15336 20154
rect 15398 20102 15410 20154
rect 15472 20102 15474 20154
rect 15312 20100 15336 20102
rect 15392 20100 15416 20102
rect 15472 20100 15496 20102
rect 15256 20080 15552 20100
rect 18256 20156 18552 20176
rect 18312 20154 18336 20156
rect 18392 20154 18416 20156
rect 18472 20154 18496 20156
rect 18334 20102 18336 20154
rect 18398 20102 18410 20154
rect 18472 20102 18474 20154
rect 18312 20100 18336 20102
rect 18392 20100 18416 20102
rect 18472 20100 18496 20102
rect 18256 20080 18552 20100
rect 21256 20156 21552 20176
rect 21312 20154 21336 20156
rect 21392 20154 21416 20156
rect 21472 20154 21496 20156
rect 21334 20102 21336 20154
rect 21398 20102 21410 20154
rect 21472 20102 21474 20154
rect 21312 20100 21336 20102
rect 21392 20100 21416 20102
rect 21472 20100 21496 20102
rect 21256 20080 21552 20100
rect 1756 19612 2052 19632
rect 1812 19610 1836 19612
rect 1892 19610 1916 19612
rect 1972 19610 1996 19612
rect 1834 19558 1836 19610
rect 1898 19558 1910 19610
rect 1972 19558 1974 19610
rect 1812 19556 1836 19558
rect 1892 19556 1916 19558
rect 1972 19556 1996 19558
rect 1756 19536 2052 19556
rect 4756 19612 5052 19632
rect 4812 19610 4836 19612
rect 4892 19610 4916 19612
rect 4972 19610 4996 19612
rect 4834 19558 4836 19610
rect 4898 19558 4910 19610
rect 4972 19558 4974 19610
rect 4812 19556 4836 19558
rect 4892 19556 4916 19558
rect 4972 19556 4996 19558
rect 4756 19536 5052 19556
rect 7756 19612 8052 19632
rect 7812 19610 7836 19612
rect 7892 19610 7916 19612
rect 7972 19610 7996 19612
rect 7834 19558 7836 19610
rect 7898 19558 7910 19610
rect 7972 19558 7974 19610
rect 7812 19556 7836 19558
rect 7892 19556 7916 19558
rect 7972 19556 7996 19558
rect 7756 19536 8052 19556
rect 10756 19612 11052 19632
rect 10812 19610 10836 19612
rect 10892 19610 10916 19612
rect 10972 19610 10996 19612
rect 10834 19558 10836 19610
rect 10898 19558 10910 19610
rect 10972 19558 10974 19610
rect 10812 19556 10836 19558
rect 10892 19556 10916 19558
rect 10972 19556 10996 19558
rect 10756 19536 11052 19556
rect 13756 19612 14052 19632
rect 13812 19610 13836 19612
rect 13892 19610 13916 19612
rect 13972 19610 13996 19612
rect 13834 19558 13836 19610
rect 13898 19558 13910 19610
rect 13972 19558 13974 19610
rect 13812 19556 13836 19558
rect 13892 19556 13916 19558
rect 13972 19556 13996 19558
rect 13756 19536 14052 19556
rect 16756 19612 17052 19632
rect 16812 19610 16836 19612
rect 16892 19610 16916 19612
rect 16972 19610 16996 19612
rect 16834 19558 16836 19610
rect 16898 19558 16910 19610
rect 16972 19558 16974 19610
rect 16812 19556 16836 19558
rect 16892 19556 16916 19558
rect 16972 19556 16996 19558
rect 16756 19536 17052 19556
rect 19756 19612 20052 19632
rect 19812 19610 19836 19612
rect 19892 19610 19916 19612
rect 19972 19610 19996 19612
rect 19834 19558 19836 19610
rect 19898 19558 19910 19610
rect 19972 19558 19974 19610
rect 19812 19556 19836 19558
rect 19892 19556 19916 19558
rect 19972 19556 19996 19558
rect 19756 19536 20052 19556
rect 22756 19612 23052 19632
rect 22812 19610 22836 19612
rect 22892 19610 22916 19612
rect 22972 19610 22996 19612
rect 22834 19558 22836 19610
rect 22898 19558 22910 19610
rect 22972 19558 22974 19610
rect 22812 19556 22836 19558
rect 22892 19556 22916 19558
rect 22972 19556 22996 19558
rect 22756 19536 23052 19556
rect 3256 19068 3552 19088
rect 3312 19066 3336 19068
rect 3392 19066 3416 19068
rect 3472 19066 3496 19068
rect 3334 19014 3336 19066
rect 3398 19014 3410 19066
rect 3472 19014 3474 19066
rect 3312 19012 3336 19014
rect 3392 19012 3416 19014
rect 3472 19012 3496 19014
rect 3256 18992 3552 19012
rect 6256 19068 6552 19088
rect 6312 19066 6336 19068
rect 6392 19066 6416 19068
rect 6472 19066 6496 19068
rect 6334 19014 6336 19066
rect 6398 19014 6410 19066
rect 6472 19014 6474 19066
rect 6312 19012 6336 19014
rect 6392 19012 6416 19014
rect 6472 19012 6496 19014
rect 6256 18992 6552 19012
rect 9256 19068 9552 19088
rect 9312 19066 9336 19068
rect 9392 19066 9416 19068
rect 9472 19066 9496 19068
rect 9334 19014 9336 19066
rect 9398 19014 9410 19066
rect 9472 19014 9474 19066
rect 9312 19012 9336 19014
rect 9392 19012 9416 19014
rect 9472 19012 9496 19014
rect 9256 18992 9552 19012
rect 12256 19068 12552 19088
rect 12312 19066 12336 19068
rect 12392 19066 12416 19068
rect 12472 19066 12496 19068
rect 12334 19014 12336 19066
rect 12398 19014 12410 19066
rect 12472 19014 12474 19066
rect 12312 19012 12336 19014
rect 12392 19012 12416 19014
rect 12472 19012 12496 19014
rect 12256 18992 12552 19012
rect 15256 19068 15552 19088
rect 15312 19066 15336 19068
rect 15392 19066 15416 19068
rect 15472 19066 15496 19068
rect 15334 19014 15336 19066
rect 15398 19014 15410 19066
rect 15472 19014 15474 19066
rect 15312 19012 15336 19014
rect 15392 19012 15416 19014
rect 15472 19012 15496 19014
rect 15256 18992 15552 19012
rect 18256 19068 18552 19088
rect 18312 19066 18336 19068
rect 18392 19066 18416 19068
rect 18472 19066 18496 19068
rect 18334 19014 18336 19066
rect 18398 19014 18410 19066
rect 18472 19014 18474 19066
rect 18312 19012 18336 19014
rect 18392 19012 18416 19014
rect 18472 19012 18496 19014
rect 18256 18992 18552 19012
rect 21256 19068 21552 19088
rect 21312 19066 21336 19068
rect 21392 19066 21416 19068
rect 21472 19066 21496 19068
rect 21334 19014 21336 19066
rect 21398 19014 21410 19066
rect 21472 19014 21474 19066
rect 21312 19012 21336 19014
rect 21392 19012 21416 19014
rect 21472 19012 21496 19014
rect 21256 18992 21552 19012
rect 1756 18524 2052 18544
rect 1812 18522 1836 18524
rect 1892 18522 1916 18524
rect 1972 18522 1996 18524
rect 1834 18470 1836 18522
rect 1898 18470 1910 18522
rect 1972 18470 1974 18522
rect 1812 18468 1836 18470
rect 1892 18468 1916 18470
rect 1972 18468 1996 18470
rect 1756 18448 2052 18468
rect 4756 18524 5052 18544
rect 4812 18522 4836 18524
rect 4892 18522 4916 18524
rect 4972 18522 4996 18524
rect 4834 18470 4836 18522
rect 4898 18470 4910 18522
rect 4972 18470 4974 18522
rect 4812 18468 4836 18470
rect 4892 18468 4916 18470
rect 4972 18468 4996 18470
rect 4756 18448 5052 18468
rect 7756 18524 8052 18544
rect 7812 18522 7836 18524
rect 7892 18522 7916 18524
rect 7972 18522 7996 18524
rect 7834 18470 7836 18522
rect 7898 18470 7910 18522
rect 7972 18470 7974 18522
rect 7812 18468 7836 18470
rect 7892 18468 7916 18470
rect 7972 18468 7996 18470
rect 7756 18448 8052 18468
rect 10756 18524 11052 18544
rect 10812 18522 10836 18524
rect 10892 18522 10916 18524
rect 10972 18522 10996 18524
rect 10834 18470 10836 18522
rect 10898 18470 10910 18522
rect 10972 18470 10974 18522
rect 10812 18468 10836 18470
rect 10892 18468 10916 18470
rect 10972 18468 10996 18470
rect 10756 18448 11052 18468
rect 13756 18524 14052 18544
rect 13812 18522 13836 18524
rect 13892 18522 13916 18524
rect 13972 18522 13996 18524
rect 13834 18470 13836 18522
rect 13898 18470 13910 18522
rect 13972 18470 13974 18522
rect 13812 18468 13836 18470
rect 13892 18468 13916 18470
rect 13972 18468 13996 18470
rect 13756 18448 14052 18468
rect 16756 18524 17052 18544
rect 16812 18522 16836 18524
rect 16892 18522 16916 18524
rect 16972 18522 16996 18524
rect 16834 18470 16836 18522
rect 16898 18470 16910 18522
rect 16972 18470 16974 18522
rect 16812 18468 16836 18470
rect 16892 18468 16916 18470
rect 16972 18468 16996 18470
rect 16756 18448 17052 18468
rect 19756 18524 20052 18544
rect 19812 18522 19836 18524
rect 19892 18522 19916 18524
rect 19972 18522 19996 18524
rect 19834 18470 19836 18522
rect 19898 18470 19910 18522
rect 19972 18470 19974 18522
rect 19812 18468 19836 18470
rect 19892 18468 19916 18470
rect 19972 18468 19996 18470
rect 19756 18448 20052 18468
rect 22756 18524 23052 18544
rect 22812 18522 22836 18524
rect 22892 18522 22916 18524
rect 22972 18522 22996 18524
rect 22834 18470 22836 18522
rect 22898 18470 22910 18522
rect 22972 18470 22974 18522
rect 22812 18468 22836 18470
rect 22892 18468 22916 18470
rect 22972 18468 22996 18470
rect 22756 18448 23052 18468
rect 3256 17980 3552 18000
rect 3312 17978 3336 17980
rect 3392 17978 3416 17980
rect 3472 17978 3496 17980
rect 3334 17926 3336 17978
rect 3398 17926 3410 17978
rect 3472 17926 3474 17978
rect 3312 17924 3336 17926
rect 3392 17924 3416 17926
rect 3472 17924 3496 17926
rect 3256 17904 3552 17924
rect 6256 17980 6552 18000
rect 6312 17978 6336 17980
rect 6392 17978 6416 17980
rect 6472 17978 6496 17980
rect 6334 17926 6336 17978
rect 6398 17926 6410 17978
rect 6472 17926 6474 17978
rect 6312 17924 6336 17926
rect 6392 17924 6416 17926
rect 6472 17924 6496 17926
rect 6256 17904 6552 17924
rect 9256 17980 9552 18000
rect 9312 17978 9336 17980
rect 9392 17978 9416 17980
rect 9472 17978 9496 17980
rect 9334 17926 9336 17978
rect 9398 17926 9410 17978
rect 9472 17926 9474 17978
rect 9312 17924 9336 17926
rect 9392 17924 9416 17926
rect 9472 17924 9496 17926
rect 9256 17904 9552 17924
rect 12256 17980 12552 18000
rect 12312 17978 12336 17980
rect 12392 17978 12416 17980
rect 12472 17978 12496 17980
rect 12334 17926 12336 17978
rect 12398 17926 12410 17978
rect 12472 17926 12474 17978
rect 12312 17924 12336 17926
rect 12392 17924 12416 17926
rect 12472 17924 12496 17926
rect 12256 17904 12552 17924
rect 15256 17980 15552 18000
rect 15312 17978 15336 17980
rect 15392 17978 15416 17980
rect 15472 17978 15496 17980
rect 15334 17926 15336 17978
rect 15398 17926 15410 17978
rect 15472 17926 15474 17978
rect 15312 17924 15336 17926
rect 15392 17924 15416 17926
rect 15472 17924 15496 17926
rect 15256 17904 15552 17924
rect 18256 17980 18552 18000
rect 18312 17978 18336 17980
rect 18392 17978 18416 17980
rect 18472 17978 18496 17980
rect 18334 17926 18336 17978
rect 18398 17926 18410 17978
rect 18472 17926 18474 17978
rect 18312 17924 18336 17926
rect 18392 17924 18416 17926
rect 18472 17924 18496 17926
rect 18256 17904 18552 17924
rect 21256 17980 21552 18000
rect 21312 17978 21336 17980
rect 21392 17978 21416 17980
rect 21472 17978 21496 17980
rect 21334 17926 21336 17978
rect 21398 17926 21410 17978
rect 21472 17926 21474 17978
rect 21312 17924 21336 17926
rect 21392 17924 21416 17926
rect 21472 17924 21496 17926
rect 21256 17904 21552 17924
rect 1756 17436 2052 17456
rect 1812 17434 1836 17436
rect 1892 17434 1916 17436
rect 1972 17434 1996 17436
rect 1834 17382 1836 17434
rect 1898 17382 1910 17434
rect 1972 17382 1974 17434
rect 1812 17380 1836 17382
rect 1892 17380 1916 17382
rect 1972 17380 1996 17382
rect 1756 17360 2052 17380
rect 4756 17436 5052 17456
rect 4812 17434 4836 17436
rect 4892 17434 4916 17436
rect 4972 17434 4996 17436
rect 4834 17382 4836 17434
rect 4898 17382 4910 17434
rect 4972 17382 4974 17434
rect 4812 17380 4836 17382
rect 4892 17380 4916 17382
rect 4972 17380 4996 17382
rect 4756 17360 5052 17380
rect 7756 17436 8052 17456
rect 7812 17434 7836 17436
rect 7892 17434 7916 17436
rect 7972 17434 7996 17436
rect 7834 17382 7836 17434
rect 7898 17382 7910 17434
rect 7972 17382 7974 17434
rect 7812 17380 7836 17382
rect 7892 17380 7916 17382
rect 7972 17380 7996 17382
rect 7756 17360 8052 17380
rect 10756 17436 11052 17456
rect 10812 17434 10836 17436
rect 10892 17434 10916 17436
rect 10972 17434 10996 17436
rect 10834 17382 10836 17434
rect 10898 17382 10910 17434
rect 10972 17382 10974 17434
rect 10812 17380 10836 17382
rect 10892 17380 10916 17382
rect 10972 17380 10996 17382
rect 10756 17360 11052 17380
rect 13756 17436 14052 17456
rect 13812 17434 13836 17436
rect 13892 17434 13916 17436
rect 13972 17434 13996 17436
rect 13834 17382 13836 17434
rect 13898 17382 13910 17434
rect 13972 17382 13974 17434
rect 13812 17380 13836 17382
rect 13892 17380 13916 17382
rect 13972 17380 13996 17382
rect 13756 17360 14052 17380
rect 16756 17436 17052 17456
rect 16812 17434 16836 17436
rect 16892 17434 16916 17436
rect 16972 17434 16996 17436
rect 16834 17382 16836 17434
rect 16898 17382 16910 17434
rect 16972 17382 16974 17434
rect 16812 17380 16836 17382
rect 16892 17380 16916 17382
rect 16972 17380 16996 17382
rect 16756 17360 17052 17380
rect 19756 17436 20052 17456
rect 19812 17434 19836 17436
rect 19892 17434 19916 17436
rect 19972 17434 19996 17436
rect 19834 17382 19836 17434
rect 19898 17382 19910 17434
rect 19972 17382 19974 17434
rect 19812 17380 19836 17382
rect 19892 17380 19916 17382
rect 19972 17380 19996 17382
rect 19756 17360 20052 17380
rect 22756 17436 23052 17456
rect 22812 17434 22836 17436
rect 22892 17434 22916 17436
rect 22972 17434 22996 17436
rect 22834 17382 22836 17434
rect 22898 17382 22910 17434
rect 22972 17382 22974 17434
rect 22812 17380 22836 17382
rect 22892 17380 22916 17382
rect 22972 17380 22996 17382
rect 22756 17360 23052 17380
rect 3256 16892 3552 16912
rect 3312 16890 3336 16892
rect 3392 16890 3416 16892
rect 3472 16890 3496 16892
rect 3334 16838 3336 16890
rect 3398 16838 3410 16890
rect 3472 16838 3474 16890
rect 3312 16836 3336 16838
rect 3392 16836 3416 16838
rect 3472 16836 3496 16838
rect 3256 16816 3552 16836
rect 6256 16892 6552 16912
rect 6312 16890 6336 16892
rect 6392 16890 6416 16892
rect 6472 16890 6496 16892
rect 6334 16838 6336 16890
rect 6398 16838 6410 16890
rect 6472 16838 6474 16890
rect 6312 16836 6336 16838
rect 6392 16836 6416 16838
rect 6472 16836 6496 16838
rect 6256 16816 6552 16836
rect 9256 16892 9552 16912
rect 9312 16890 9336 16892
rect 9392 16890 9416 16892
rect 9472 16890 9496 16892
rect 9334 16838 9336 16890
rect 9398 16838 9410 16890
rect 9472 16838 9474 16890
rect 9312 16836 9336 16838
rect 9392 16836 9416 16838
rect 9472 16836 9496 16838
rect 9256 16816 9552 16836
rect 12256 16892 12552 16912
rect 12312 16890 12336 16892
rect 12392 16890 12416 16892
rect 12472 16890 12496 16892
rect 12334 16838 12336 16890
rect 12398 16838 12410 16890
rect 12472 16838 12474 16890
rect 12312 16836 12336 16838
rect 12392 16836 12416 16838
rect 12472 16836 12496 16838
rect 12256 16816 12552 16836
rect 15256 16892 15552 16912
rect 15312 16890 15336 16892
rect 15392 16890 15416 16892
rect 15472 16890 15496 16892
rect 15334 16838 15336 16890
rect 15398 16838 15410 16890
rect 15472 16838 15474 16890
rect 15312 16836 15336 16838
rect 15392 16836 15416 16838
rect 15472 16836 15496 16838
rect 15256 16816 15552 16836
rect 18256 16892 18552 16912
rect 18312 16890 18336 16892
rect 18392 16890 18416 16892
rect 18472 16890 18496 16892
rect 18334 16838 18336 16890
rect 18398 16838 18410 16890
rect 18472 16838 18474 16890
rect 18312 16836 18336 16838
rect 18392 16836 18416 16838
rect 18472 16836 18496 16838
rect 18256 16816 18552 16836
rect 21256 16892 21552 16912
rect 21312 16890 21336 16892
rect 21392 16890 21416 16892
rect 21472 16890 21496 16892
rect 21334 16838 21336 16890
rect 21398 16838 21410 16890
rect 21472 16838 21474 16890
rect 21312 16836 21336 16838
rect 21392 16836 21416 16838
rect 21472 16836 21496 16838
rect 21256 16816 21552 16836
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 1756 16348 2052 16368
rect 1812 16346 1836 16348
rect 1892 16346 1916 16348
rect 1972 16346 1996 16348
rect 1834 16294 1836 16346
rect 1898 16294 1910 16346
rect 1972 16294 1974 16346
rect 1812 16292 1836 16294
rect 1892 16292 1916 16294
rect 1972 16292 1996 16294
rect 1756 16272 2052 16292
rect 4756 16348 5052 16368
rect 4812 16346 4836 16348
rect 4892 16346 4916 16348
rect 4972 16346 4996 16348
rect 4834 16294 4836 16346
rect 4898 16294 4910 16346
rect 4972 16294 4974 16346
rect 4812 16292 4836 16294
rect 4892 16292 4916 16294
rect 4972 16292 4996 16294
rect 4756 16272 5052 16292
rect 7756 16348 8052 16368
rect 7812 16346 7836 16348
rect 7892 16346 7916 16348
rect 7972 16346 7996 16348
rect 7834 16294 7836 16346
rect 7898 16294 7910 16346
rect 7972 16294 7974 16346
rect 7812 16292 7836 16294
rect 7892 16292 7916 16294
rect 7972 16292 7996 16294
rect 7756 16272 8052 16292
rect 10756 16348 11052 16368
rect 10812 16346 10836 16348
rect 10892 16346 10916 16348
rect 10972 16346 10996 16348
rect 10834 16294 10836 16346
rect 10898 16294 10910 16346
rect 10972 16294 10974 16346
rect 10812 16292 10836 16294
rect 10892 16292 10916 16294
rect 10972 16292 10996 16294
rect 10756 16272 11052 16292
rect 13756 16348 14052 16368
rect 13812 16346 13836 16348
rect 13892 16346 13916 16348
rect 13972 16346 13996 16348
rect 13834 16294 13836 16346
rect 13898 16294 13910 16346
rect 13972 16294 13974 16346
rect 13812 16292 13836 16294
rect 13892 16292 13916 16294
rect 13972 16292 13996 16294
rect 13756 16272 14052 16292
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 3256 15804 3552 15824
rect 3312 15802 3336 15804
rect 3392 15802 3416 15804
rect 3472 15802 3496 15804
rect 3334 15750 3336 15802
rect 3398 15750 3410 15802
rect 3472 15750 3474 15802
rect 3312 15748 3336 15750
rect 3392 15748 3416 15750
rect 3472 15748 3496 15750
rect 3256 15728 3552 15748
rect 6256 15804 6552 15824
rect 6312 15802 6336 15804
rect 6392 15802 6416 15804
rect 6472 15802 6496 15804
rect 6334 15750 6336 15802
rect 6398 15750 6410 15802
rect 6472 15750 6474 15802
rect 6312 15748 6336 15750
rect 6392 15748 6416 15750
rect 6472 15748 6496 15750
rect 6256 15728 6552 15748
rect 9256 15804 9552 15824
rect 9312 15802 9336 15804
rect 9392 15802 9416 15804
rect 9472 15802 9496 15804
rect 9334 15750 9336 15802
rect 9398 15750 9410 15802
rect 9472 15750 9474 15802
rect 9312 15748 9336 15750
rect 9392 15748 9416 15750
rect 9472 15748 9496 15750
rect 9256 15728 9552 15748
rect 12256 15804 12552 15824
rect 12312 15802 12336 15804
rect 12392 15802 12416 15804
rect 12472 15802 12496 15804
rect 12334 15750 12336 15802
rect 12398 15750 12410 15802
rect 12472 15750 12474 15802
rect 12312 15748 12336 15750
rect 12392 15748 12416 15750
rect 12472 15748 12496 15750
rect 12256 15728 12552 15748
rect 13832 15570 13860 15846
rect 14292 15570 14320 16526
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 16250 14412 16390
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14752 16182 14780 16662
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 14648 16176 14700 16182
rect 14648 16118 14700 16124
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 1756 15260 2052 15280
rect 1812 15258 1836 15260
rect 1892 15258 1916 15260
rect 1972 15258 1996 15260
rect 1834 15206 1836 15258
rect 1898 15206 1910 15258
rect 1972 15206 1974 15258
rect 1812 15204 1836 15206
rect 1892 15204 1916 15206
rect 1972 15204 1996 15206
rect 1756 15184 2052 15204
rect 4756 15260 5052 15280
rect 4812 15258 4836 15260
rect 4892 15258 4916 15260
rect 4972 15258 4996 15260
rect 4834 15206 4836 15258
rect 4898 15206 4910 15258
rect 4972 15206 4974 15258
rect 4812 15204 4836 15206
rect 4892 15204 4916 15206
rect 4972 15204 4996 15206
rect 4756 15184 5052 15204
rect 7756 15260 8052 15280
rect 7812 15258 7836 15260
rect 7892 15258 7916 15260
rect 7972 15258 7996 15260
rect 7834 15206 7836 15258
rect 7898 15206 7910 15258
rect 7972 15206 7974 15258
rect 7812 15204 7836 15206
rect 7892 15204 7916 15206
rect 7972 15204 7996 15206
rect 7756 15184 8052 15204
rect 10756 15260 11052 15280
rect 10812 15258 10836 15260
rect 10892 15258 10916 15260
rect 10972 15258 10996 15260
rect 10834 15206 10836 15258
rect 10898 15206 10910 15258
rect 10972 15206 10974 15258
rect 10812 15204 10836 15206
rect 10892 15204 10916 15206
rect 10972 15204 10996 15206
rect 10756 15184 11052 15204
rect 12820 15162 12848 15438
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 3256 14716 3552 14736
rect 3312 14714 3336 14716
rect 3392 14714 3416 14716
rect 3472 14714 3496 14716
rect 3334 14662 3336 14714
rect 3398 14662 3410 14714
rect 3472 14662 3474 14714
rect 3312 14660 3336 14662
rect 3392 14660 3416 14662
rect 3472 14660 3496 14662
rect 3256 14640 3552 14660
rect 6256 14716 6552 14736
rect 6312 14714 6336 14716
rect 6392 14714 6416 14716
rect 6472 14714 6496 14716
rect 6334 14662 6336 14714
rect 6398 14662 6410 14714
rect 6472 14662 6474 14714
rect 6312 14660 6336 14662
rect 6392 14660 6416 14662
rect 6472 14660 6496 14662
rect 6256 14640 6552 14660
rect 9256 14716 9552 14736
rect 9312 14714 9336 14716
rect 9392 14714 9416 14716
rect 9472 14714 9496 14716
rect 9334 14662 9336 14714
rect 9398 14662 9410 14714
rect 9472 14662 9474 14714
rect 9312 14660 9336 14662
rect 9392 14660 9416 14662
rect 9472 14660 9496 14662
rect 9256 14640 9552 14660
rect 12256 14716 12552 14736
rect 12312 14714 12336 14716
rect 12392 14714 12416 14716
rect 12472 14714 12496 14716
rect 12334 14662 12336 14714
rect 12398 14662 12410 14714
rect 12472 14662 12474 14714
rect 12312 14660 12336 14662
rect 12392 14660 12416 14662
rect 12472 14660 12496 14662
rect 12256 14640 12552 14660
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 1756 14172 2052 14192
rect 1812 14170 1836 14172
rect 1892 14170 1916 14172
rect 1972 14170 1996 14172
rect 1834 14118 1836 14170
rect 1898 14118 1910 14170
rect 1972 14118 1974 14170
rect 1812 14116 1836 14118
rect 1892 14116 1916 14118
rect 1972 14116 1996 14118
rect 1756 14096 2052 14116
rect 4756 14172 5052 14192
rect 4812 14170 4836 14172
rect 4892 14170 4916 14172
rect 4972 14170 4996 14172
rect 4834 14118 4836 14170
rect 4898 14118 4910 14170
rect 4972 14118 4974 14170
rect 4812 14116 4836 14118
rect 4892 14116 4916 14118
rect 4972 14116 4996 14118
rect 4756 14096 5052 14116
rect 7756 14172 8052 14192
rect 7812 14170 7836 14172
rect 7892 14170 7916 14172
rect 7972 14170 7996 14172
rect 7834 14118 7836 14170
rect 7898 14118 7910 14170
rect 7972 14118 7974 14170
rect 7812 14116 7836 14118
rect 7892 14116 7916 14118
rect 7972 14116 7996 14118
rect 7756 14096 8052 14116
rect 10756 14172 11052 14192
rect 10812 14170 10836 14172
rect 10892 14170 10916 14172
rect 10972 14170 10996 14172
rect 10834 14118 10836 14170
rect 10898 14118 10910 14170
rect 10972 14118 10974 14170
rect 10812 14116 10836 14118
rect 10892 14116 10916 14118
rect 10972 14116 10996 14118
rect 10756 14096 11052 14116
rect 8482 13968 8538 13977
rect 8482 13903 8484 13912
rect 8536 13903 8538 13912
rect 8484 13874 8536 13880
rect 110 13696 166 13705
rect 110 13631 166 13640
rect 124 12753 152 13631
rect 3256 13628 3552 13648
rect 3312 13626 3336 13628
rect 3392 13626 3416 13628
rect 3472 13626 3496 13628
rect 3334 13574 3336 13626
rect 3398 13574 3410 13626
rect 3472 13574 3474 13626
rect 3312 13572 3336 13574
rect 3392 13572 3416 13574
rect 3472 13572 3496 13574
rect 3256 13552 3552 13572
rect 6256 13628 6552 13648
rect 6312 13626 6336 13628
rect 6392 13626 6416 13628
rect 6472 13626 6496 13628
rect 6334 13574 6336 13626
rect 6398 13574 6410 13626
rect 6472 13574 6474 13626
rect 6312 13572 6336 13574
rect 6392 13572 6416 13574
rect 6472 13572 6496 13574
rect 6256 13552 6552 13572
rect 8496 13190 8524 13874
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 1756 13084 2052 13104
rect 1812 13082 1836 13084
rect 1892 13082 1916 13084
rect 1972 13082 1996 13084
rect 1834 13030 1836 13082
rect 1898 13030 1910 13082
rect 1972 13030 1974 13082
rect 1812 13028 1836 13030
rect 1892 13028 1916 13030
rect 1972 13028 1996 13030
rect 1756 13008 2052 13028
rect 4756 13084 5052 13104
rect 4812 13082 4836 13084
rect 4892 13082 4916 13084
rect 4972 13082 4996 13084
rect 4834 13030 4836 13082
rect 4898 13030 4910 13082
rect 4972 13030 4974 13082
rect 4812 13028 4836 13030
rect 4892 13028 4916 13030
rect 4972 13028 4996 13030
rect 4756 13008 5052 13028
rect 7756 13084 8052 13104
rect 7812 13082 7836 13084
rect 7892 13082 7916 13084
rect 7972 13082 7996 13084
rect 7834 13030 7836 13082
rect 7898 13030 7910 13082
rect 7972 13030 7974 13082
rect 7812 13028 7836 13030
rect 7892 13028 7916 13030
rect 7972 13028 7996 13030
rect 7756 13008 8052 13028
rect 110 12744 166 12753
rect 110 12679 166 12688
rect 3256 12540 3552 12560
rect 3312 12538 3336 12540
rect 3392 12538 3416 12540
rect 3472 12538 3496 12540
rect 3334 12486 3336 12538
rect 3398 12486 3410 12538
rect 3472 12486 3474 12538
rect 3312 12484 3336 12486
rect 3392 12484 3416 12486
rect 3472 12484 3496 12486
rect 3256 12464 3552 12484
rect 6256 12540 6552 12560
rect 6312 12538 6336 12540
rect 6392 12538 6416 12540
rect 6472 12538 6496 12540
rect 6334 12486 6336 12538
rect 6398 12486 6410 12538
rect 6472 12486 6474 12538
rect 6312 12484 6336 12486
rect 6392 12484 6416 12486
rect 6472 12484 6496 12486
rect 6256 12464 6552 12484
rect 1756 11996 2052 12016
rect 1812 11994 1836 11996
rect 1892 11994 1916 11996
rect 1972 11994 1996 11996
rect 1834 11942 1836 11994
rect 1898 11942 1910 11994
rect 1972 11942 1974 11994
rect 1812 11940 1836 11942
rect 1892 11940 1916 11942
rect 1972 11940 1996 11942
rect 1756 11920 2052 11940
rect 4756 11996 5052 12016
rect 4812 11994 4836 11996
rect 4892 11994 4916 11996
rect 4972 11994 4996 11996
rect 4834 11942 4836 11994
rect 4898 11942 4910 11994
rect 4972 11942 4974 11994
rect 4812 11940 4836 11942
rect 4892 11940 4916 11942
rect 4972 11940 4996 11942
rect 4756 11920 5052 11940
rect 7756 11996 8052 12016
rect 7812 11994 7836 11996
rect 7892 11994 7916 11996
rect 7972 11994 7996 11996
rect 7834 11942 7836 11994
rect 7898 11942 7910 11994
rect 7972 11942 7974 11994
rect 7812 11940 7836 11942
rect 7892 11940 7916 11942
rect 7972 11940 7996 11942
rect 7756 11920 8052 11940
rect 3256 11452 3552 11472
rect 3312 11450 3336 11452
rect 3392 11450 3416 11452
rect 3472 11450 3496 11452
rect 3334 11398 3336 11450
rect 3398 11398 3410 11450
rect 3472 11398 3474 11450
rect 3312 11396 3336 11398
rect 3392 11396 3416 11398
rect 3472 11396 3496 11398
rect 3256 11376 3552 11396
rect 6256 11452 6552 11472
rect 6312 11450 6336 11452
rect 6392 11450 6416 11452
rect 6472 11450 6496 11452
rect 6334 11398 6336 11450
rect 6398 11398 6410 11450
rect 6472 11398 6474 11450
rect 6312 11396 6336 11398
rect 6392 11396 6416 11398
rect 6472 11396 6496 11398
rect 6256 11376 6552 11396
rect 1756 10908 2052 10928
rect 1812 10906 1836 10908
rect 1892 10906 1916 10908
rect 1972 10906 1996 10908
rect 1834 10854 1836 10906
rect 1898 10854 1910 10906
rect 1972 10854 1974 10906
rect 1812 10852 1836 10854
rect 1892 10852 1916 10854
rect 1972 10852 1996 10854
rect 1756 10832 2052 10852
rect 4756 10908 5052 10928
rect 4812 10906 4836 10908
rect 4892 10906 4916 10908
rect 4972 10906 4996 10908
rect 4834 10854 4836 10906
rect 4898 10854 4910 10906
rect 4972 10854 4974 10906
rect 4812 10852 4836 10854
rect 4892 10852 4916 10854
rect 4972 10852 4996 10854
rect 4756 10832 5052 10852
rect 7756 10908 8052 10928
rect 7812 10906 7836 10908
rect 7892 10906 7916 10908
rect 7972 10906 7996 10908
rect 7834 10854 7836 10906
rect 7898 10854 7910 10906
rect 7972 10854 7974 10906
rect 7812 10852 7836 10854
rect 7892 10852 7916 10854
rect 7972 10852 7996 10854
rect 7756 10832 8052 10852
rect 3256 10364 3552 10384
rect 3312 10362 3336 10364
rect 3392 10362 3416 10364
rect 3472 10362 3496 10364
rect 3334 10310 3336 10362
rect 3398 10310 3410 10362
rect 3472 10310 3474 10362
rect 3312 10308 3336 10310
rect 3392 10308 3416 10310
rect 3472 10308 3496 10310
rect 3256 10288 3552 10308
rect 6256 10364 6552 10384
rect 6312 10362 6336 10364
rect 6392 10362 6416 10364
rect 6472 10362 6496 10364
rect 6334 10310 6336 10362
rect 6398 10310 6410 10362
rect 6472 10310 6474 10362
rect 6312 10308 6336 10310
rect 6392 10308 6416 10310
rect 6472 10308 6496 10310
rect 6256 10288 6552 10308
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 1756 9820 2052 9840
rect 1812 9818 1836 9820
rect 1892 9818 1916 9820
rect 1972 9818 1996 9820
rect 1834 9766 1836 9818
rect 1898 9766 1910 9818
rect 1972 9766 1974 9818
rect 1812 9764 1836 9766
rect 1892 9764 1916 9766
rect 1972 9764 1996 9766
rect 1756 9744 2052 9764
rect 4756 9820 5052 9840
rect 4812 9818 4836 9820
rect 4892 9818 4916 9820
rect 4972 9818 4996 9820
rect 4834 9766 4836 9818
rect 4898 9766 4910 9818
rect 4972 9766 4974 9818
rect 4812 9764 4836 9766
rect 4892 9764 4916 9766
rect 4972 9764 4996 9766
rect 4756 9744 5052 9764
rect 7024 9722 7052 9930
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7116 9382 7144 10066
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7484 9450 7512 9930
rect 7756 9820 8052 9840
rect 7812 9818 7836 9820
rect 7892 9818 7916 9820
rect 7972 9818 7996 9820
rect 7834 9766 7836 9818
rect 7898 9766 7910 9818
rect 7972 9766 7974 9818
rect 7812 9764 7836 9766
rect 7892 9764 7916 9766
rect 7972 9764 7996 9766
rect 7756 9744 8052 9764
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 3256 9276 3552 9296
rect 3312 9274 3336 9276
rect 3392 9274 3416 9276
rect 3472 9274 3496 9276
rect 3334 9222 3336 9274
rect 3398 9222 3410 9274
rect 3472 9222 3474 9274
rect 3312 9220 3336 9222
rect 3392 9220 3416 9222
rect 3472 9220 3496 9222
rect 3256 9200 3552 9220
rect 6256 9276 6552 9296
rect 6312 9274 6336 9276
rect 6392 9274 6416 9276
rect 6472 9274 6496 9276
rect 6334 9222 6336 9274
rect 6398 9222 6410 9274
rect 6472 9222 6474 9274
rect 6312 9220 6336 9222
rect 6392 9220 6416 9222
rect 6472 9220 6496 9222
rect 6256 9200 6552 9220
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 1756 8732 2052 8752
rect 1812 8730 1836 8732
rect 1892 8730 1916 8732
rect 1972 8730 1996 8732
rect 1834 8678 1836 8730
rect 1898 8678 1910 8730
rect 1972 8678 1974 8730
rect 1812 8676 1836 8678
rect 1892 8676 1916 8678
rect 1972 8676 1996 8678
rect 1756 8656 2052 8676
rect 4756 8732 5052 8752
rect 4812 8730 4836 8732
rect 4892 8730 4916 8732
rect 4972 8730 4996 8732
rect 4834 8678 4836 8730
rect 4898 8678 4910 8730
rect 4972 8678 4974 8730
rect 4812 8676 4836 8678
rect 4892 8676 4916 8678
rect 4972 8676 4996 8678
rect 4756 8656 5052 8676
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 3256 8188 3552 8208
rect 3312 8186 3336 8188
rect 3392 8186 3416 8188
rect 3472 8186 3496 8188
rect 3334 8134 3336 8186
rect 3398 8134 3410 8186
rect 3472 8134 3474 8186
rect 3312 8132 3336 8134
rect 3392 8132 3416 8134
rect 3472 8132 3496 8134
rect 3256 8112 3552 8132
rect 1756 7644 2052 7664
rect 1812 7642 1836 7644
rect 1892 7642 1916 7644
rect 1972 7642 1996 7644
rect 1834 7590 1836 7642
rect 1898 7590 1910 7642
rect 1972 7590 1974 7642
rect 1812 7588 1836 7590
rect 1892 7588 1916 7590
rect 1972 7588 1996 7590
rect 1756 7568 2052 7588
rect 4756 7644 5052 7664
rect 4812 7642 4836 7644
rect 4892 7642 4916 7644
rect 4972 7642 4996 7644
rect 4834 7590 4836 7642
rect 4898 7590 4910 7642
rect 4972 7590 4974 7642
rect 4812 7588 4836 7590
rect 4892 7588 4916 7590
rect 4972 7588 4996 7590
rect 4756 7568 5052 7588
rect 3256 7100 3552 7120
rect 3312 7098 3336 7100
rect 3392 7098 3416 7100
rect 3472 7098 3496 7100
rect 3334 7046 3336 7098
rect 3398 7046 3410 7098
rect 3472 7046 3474 7098
rect 3312 7044 3336 7046
rect 3392 7044 3416 7046
rect 3472 7044 3496 7046
rect 3256 7024 3552 7044
rect 1756 6556 2052 6576
rect 1812 6554 1836 6556
rect 1892 6554 1916 6556
rect 1972 6554 1996 6556
rect 1834 6502 1836 6554
rect 1898 6502 1910 6554
rect 1972 6502 1974 6554
rect 1812 6500 1836 6502
rect 1892 6500 1916 6502
rect 1972 6500 1996 6502
rect 1756 6480 2052 6500
rect 4756 6556 5052 6576
rect 4812 6554 4836 6556
rect 4892 6554 4916 6556
rect 4972 6554 4996 6556
rect 4834 6502 4836 6554
rect 4898 6502 4910 6554
rect 4972 6502 4974 6554
rect 4812 6500 4836 6502
rect 4892 6500 4916 6502
rect 4972 6500 4996 6502
rect 4756 6480 5052 6500
rect 5736 6322 5764 8230
rect 6196 7954 6224 8774
rect 6256 8188 6552 8208
rect 6312 8186 6336 8188
rect 6392 8186 6416 8188
rect 6472 8186 6496 8188
rect 6334 8134 6336 8186
rect 6398 8134 6410 8186
rect 6472 8134 6474 8186
rect 6312 8132 6336 8134
rect 6392 8132 6416 8134
rect 6472 8132 6496 8134
rect 6256 8112 6552 8132
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6256 7100 6552 7120
rect 6312 7098 6336 7100
rect 6392 7098 6416 7100
rect 6472 7098 6496 7100
rect 6334 7046 6336 7098
rect 6398 7046 6410 7098
rect 6472 7046 6474 7098
rect 6312 7044 6336 7046
rect 6392 7044 6416 7046
rect 6472 7044 6496 7046
rect 6256 7024 6552 7044
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 3256 6012 3552 6032
rect 3312 6010 3336 6012
rect 3392 6010 3416 6012
rect 3472 6010 3496 6012
rect 3334 5958 3336 6010
rect 3398 5958 3410 6010
rect 3472 5958 3474 6010
rect 3312 5956 3336 5958
rect 3392 5956 3416 5958
rect 3472 5956 3496 5958
rect 3256 5936 3552 5956
rect 5736 5914 5764 6258
rect 6256 6012 6552 6032
rect 6312 6010 6336 6012
rect 6392 6010 6416 6012
rect 6472 6010 6496 6012
rect 6334 5958 6336 6010
rect 6398 5958 6410 6010
rect 6472 5958 6474 6010
rect 6312 5956 6336 5958
rect 6392 5956 6416 5958
rect 6472 5956 6496 5958
rect 6256 5936 6552 5956
rect 6748 5914 6776 6734
rect 7116 6254 7144 9318
rect 7484 9178 7512 9386
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7208 8294 7236 8910
rect 7756 8732 8052 8752
rect 7812 8730 7836 8732
rect 7892 8730 7916 8732
rect 7972 8730 7996 8732
rect 7834 8678 7836 8730
rect 7898 8678 7910 8730
rect 7972 8678 7974 8730
rect 7812 8676 7836 8678
rect 7892 8676 7916 8678
rect 7972 8676 7996 8678
rect 7756 8656 8052 8676
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7208 8022 7236 8230
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7944 7886 7972 8230
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7484 7410 7512 7754
rect 7756 7644 8052 7664
rect 7812 7642 7836 7644
rect 7892 7642 7916 7644
rect 7972 7642 7996 7644
rect 7834 7590 7836 7642
rect 7898 7590 7910 7642
rect 7972 7590 7974 7642
rect 7812 7588 7836 7590
rect 7892 7588 7916 7590
rect 7972 7588 7996 7590
rect 7756 7568 8052 7588
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7116 5574 7144 6190
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 1756 5468 2052 5488
rect 1812 5466 1836 5468
rect 1892 5466 1916 5468
rect 1972 5466 1996 5468
rect 1834 5414 1836 5466
rect 1898 5414 1910 5466
rect 1972 5414 1974 5466
rect 1812 5412 1836 5414
rect 1892 5412 1916 5414
rect 1972 5412 1996 5414
rect 1756 5392 2052 5412
rect 4756 5468 5052 5488
rect 4812 5466 4836 5468
rect 4892 5466 4916 5468
rect 4972 5466 4996 5468
rect 4834 5414 4836 5466
rect 4898 5414 4910 5466
rect 4972 5414 4974 5466
rect 4812 5412 4836 5414
rect 4892 5412 4916 5414
rect 4972 5412 4996 5414
rect 4756 5392 5052 5412
rect 7208 5370 7236 6394
rect 7392 6254 7420 6666
rect 7484 6644 7512 7346
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6798 7604 7142
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7564 6656 7616 6662
rect 7484 6616 7564 6644
rect 7564 6598 7616 6604
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5914 7420 6190
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7576 5624 7604 6598
rect 7668 5914 7696 6802
rect 8128 6798 8156 13126
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 12306 8708 12718
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8220 11898 8248 12242
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8312 11898 8340 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8312 10810 8340 11834
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8588 11014 8616 11562
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8220 9586 8248 10542
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8220 9110 8248 9522
rect 8312 9178 8340 10746
rect 8588 10588 8616 10950
rect 8680 10742 8708 12242
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8668 10600 8720 10606
rect 8588 10560 8668 10588
rect 8668 10542 8720 10548
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8588 9586 8616 10406
rect 8680 9976 8708 10542
rect 8772 10266 8800 10610
rect 8864 10470 8892 13670
rect 9256 13628 9552 13648
rect 9312 13626 9336 13628
rect 9392 13626 9416 13628
rect 9472 13626 9496 13628
rect 9334 13574 9336 13626
rect 9398 13574 9410 13626
rect 9472 13574 9474 13626
rect 9312 13572 9336 13574
rect 9392 13572 9416 13574
rect 9472 13572 9496 13574
rect 9256 13552 9552 13572
rect 10756 13084 11052 13104
rect 10812 13082 10836 13084
rect 10892 13082 10916 13084
rect 10972 13082 10996 13084
rect 10834 13030 10836 13082
rect 10898 13030 10910 13082
rect 10972 13030 10974 13082
rect 10812 13028 10836 13030
rect 10892 13028 10916 13030
rect 10972 13028 10996 13030
rect 10756 13008 11052 13028
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9140 12442 9168 12786
rect 9256 12540 9552 12560
rect 9312 12538 9336 12540
rect 9392 12538 9416 12540
rect 9472 12538 9496 12540
rect 9334 12486 9336 12538
rect 9398 12486 9410 12538
rect 9472 12486 9474 12538
rect 9312 12484 9336 12486
rect 9392 12484 9416 12486
rect 9472 12484 9496 12486
rect 9256 12464 9552 12484
rect 9128 12436 9180 12442
rect 8956 12396 9128 12424
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8760 9988 8812 9994
rect 8680 9948 8760 9976
rect 8760 9930 8812 9936
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8220 8634 8248 8910
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8294 8340 8910
rect 8588 8906 8616 9522
rect 8772 9450 8800 9930
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8956 8498 8984 12396
rect 9128 12378 9180 12384
rect 11440 12238 11468 14214
rect 11532 13734 11560 14350
rect 12636 14278 12664 14894
rect 12912 14482 12940 14894
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11532 13530 11560 13670
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11532 12986 11560 13466
rect 11716 13190 11744 13670
rect 12256 13628 12552 13648
rect 12312 13626 12336 13628
rect 12392 13626 12416 13628
rect 12472 13626 12496 13628
rect 12334 13574 12336 13626
rect 12398 13574 12410 13626
rect 12472 13574 12474 13626
rect 12312 13572 12336 13574
rect 12392 13572 12416 13574
rect 12472 13572 12496 13574
rect 12256 13552 12552 13572
rect 12728 13530 12756 14282
rect 13004 14074 13032 15302
rect 13372 15094 13400 15302
rect 13756 15260 14052 15280
rect 13812 15258 13836 15260
rect 13892 15258 13916 15260
rect 13972 15258 13996 15260
rect 13834 15206 13836 15258
rect 13898 15206 13910 15258
rect 13972 15206 13974 15258
rect 13812 15204 13836 15206
rect 13892 15204 13916 15206
rect 13972 15204 13996 15206
rect 13756 15184 14052 15204
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 13280 12986 13308 14010
rect 13372 14006 13400 14350
rect 13360 14000 13412 14006
rect 13360 13942 13412 13948
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13464 13394 13492 13874
rect 13556 13870 13584 14350
rect 13648 14074 13676 14350
rect 13756 14172 14052 14192
rect 13812 14170 13836 14172
rect 13892 14170 13916 14172
rect 13972 14170 13996 14172
rect 13834 14118 13836 14170
rect 13898 14118 13910 14170
rect 13972 14118 13974 14170
rect 13812 14116 13836 14118
rect 13892 14116 13916 14118
rect 13972 14116 13996 14118
rect 13756 14096 14052 14116
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 14108 13977 14136 14554
rect 14200 14482 14228 14962
rect 14292 14521 14320 15506
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 14618 14596 15438
rect 14660 15366 14688 16118
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 15162 14688 15302
rect 14752 15162 14780 16118
rect 16132 16046 16160 16390
rect 16316 16250 16344 16526
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15256 15804 15552 15824
rect 15312 15802 15336 15804
rect 15392 15802 15416 15804
rect 15472 15802 15496 15804
rect 15334 15750 15336 15802
rect 15398 15750 15410 15802
rect 15472 15750 15474 15802
rect 15312 15748 15336 15750
rect 15392 15748 15416 15750
rect 15472 15748 15496 15750
rect 15256 15728 15552 15748
rect 16132 15502 16160 15982
rect 16500 15706 16528 16526
rect 16756 16348 17052 16368
rect 16812 16346 16836 16348
rect 16892 16346 16916 16348
rect 16972 16346 16996 16348
rect 16834 16294 16836 16346
rect 16898 16294 16910 16346
rect 16972 16294 16974 16346
rect 16812 16292 16836 16294
rect 16892 16292 16916 16294
rect 16972 16292 16996 16294
rect 16756 16272 17052 16292
rect 17144 15910 17172 16526
rect 19756 16348 20052 16368
rect 19812 16346 19836 16348
rect 19892 16346 19916 16348
rect 19972 16346 19996 16348
rect 19834 16294 19836 16346
rect 19898 16294 19910 16346
rect 19972 16294 19974 16346
rect 19812 16292 19836 16294
rect 19892 16292 19916 16294
rect 19972 16292 19996 16294
rect 19756 16272 20052 16292
rect 22756 16348 23052 16368
rect 22812 16346 22836 16348
rect 22892 16346 22916 16348
rect 22972 16346 22996 16348
rect 22834 16294 22836 16346
rect 22898 16294 22910 16346
rect 22972 16294 22974 16346
rect 22812 16292 22836 16294
rect 22892 16292 22916 16294
rect 22972 16292 22996 16294
rect 22756 16272 23052 16292
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 17144 15570 17172 15846
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15256 14716 15552 14736
rect 15312 14714 15336 14716
rect 15392 14714 15416 14716
rect 15472 14714 15496 14716
rect 15334 14662 15336 14714
rect 15398 14662 15410 14714
rect 15472 14662 15474 14714
rect 15312 14660 15336 14662
rect 15392 14660 15416 14662
rect 15472 14660 15496 14662
rect 15256 14640 15552 14660
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14278 14512 14334 14521
rect 14188 14476 14240 14482
rect 15672 14482 15700 14758
rect 14278 14447 14334 14456
rect 14372 14476 14424 14482
rect 14188 14418 14240 14424
rect 14372 14418 14424 14424
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 14094 13968 14150 13977
rect 14384 13938 14412 14418
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 14074 15516 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 14094 13903 14150 13912
rect 14372 13932 14424 13938
rect 13544 13864 13596 13870
rect 14108 13814 14136 13903
rect 14372 13874 14424 13880
rect 13544 13806 13596 13812
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 11532 12442 11560 12922
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11808 12306 11836 12718
rect 12256 12540 12552 12560
rect 12312 12538 12336 12540
rect 12392 12538 12416 12540
rect 12472 12538 12496 12540
rect 12334 12486 12336 12538
rect 12398 12486 12410 12538
rect 12472 12486 12474 12538
rect 12312 12484 12336 12486
rect 12392 12484 12416 12486
rect 12472 12484 12496 12486
rect 12256 12464 12552 12484
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9048 10198 9076 10678
rect 9036 10192 9088 10198
rect 9036 10134 9088 10140
rect 9140 9518 9168 11630
rect 9256 11452 9552 11472
rect 9312 11450 9336 11452
rect 9392 11450 9416 11452
rect 9472 11450 9496 11452
rect 9334 11398 9336 11450
rect 9398 11398 9410 11450
rect 9472 11398 9474 11450
rect 9312 11396 9336 11398
rect 9392 11396 9416 11398
rect 9472 11396 9496 11398
rect 9256 11376 9552 11396
rect 9600 11286 9628 11630
rect 9784 11354 9812 11698
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9256 10364 9552 10384
rect 9312 10362 9336 10364
rect 9392 10362 9416 10364
rect 9472 10362 9496 10364
rect 9334 10310 9336 10362
rect 9398 10310 9410 10362
rect 9472 10310 9474 10362
rect 9312 10308 9336 10310
rect 9392 10308 9416 10310
rect 9472 10308 9496 10310
rect 9256 10288 9552 10308
rect 9784 9586 9812 11290
rect 9876 10062 9904 12106
rect 10756 11996 11052 12016
rect 10812 11994 10836 11996
rect 10892 11994 10916 11996
rect 10972 11994 10996 11996
rect 10834 11942 10836 11994
rect 10898 11942 10910 11994
rect 10972 11942 10974 11994
rect 10812 11940 10836 11942
rect 10892 11940 10916 11942
rect 10972 11940 10996 11942
rect 10756 11920 11052 11940
rect 11440 11558 11468 12174
rect 11808 11830 11836 12242
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12268 11898 12296 12106
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10336 10266 10364 10610
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 9722 9904 9998
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9048 9178 9076 9454
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9048 8566 9076 9114
rect 9140 9042 9168 9454
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9256 9276 9552 9296
rect 9312 9274 9336 9276
rect 9392 9274 9416 9276
rect 9472 9274 9496 9276
rect 9334 9222 9336 9274
rect 9398 9222 9410 9274
rect 9472 9222 9474 9274
rect 9312 9220 9336 9222
rect 9392 9220 9416 9222
rect 9472 9220 9496 9222
rect 9256 9200 9552 9220
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8956 8090 8984 8434
rect 9876 8294 9904 8842
rect 9968 8498 9996 9318
rect 10428 9042 10456 10950
rect 10756 10908 11052 10928
rect 10812 10906 10836 10908
rect 10892 10906 10916 10908
rect 10972 10906 10996 10908
rect 10834 10854 10836 10906
rect 10898 10854 10910 10906
rect 10972 10854 10974 10906
rect 10812 10852 10836 10854
rect 10892 10852 10916 10854
rect 10972 10852 10996 10854
rect 10756 10832 11052 10852
rect 11164 10130 11192 11018
rect 11348 10742 11376 11154
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9586 10640 9862
rect 10756 9820 11052 9840
rect 10812 9818 10836 9820
rect 10892 9818 10916 9820
rect 10972 9818 10996 9820
rect 10834 9766 10836 9818
rect 10898 9766 10910 9818
rect 10972 9766 10974 9818
rect 10812 9764 10836 9766
rect 10892 9764 10916 9766
rect 10972 9764 10996 9766
rect 10756 9744 11052 9764
rect 11164 9722 11192 10066
rect 11440 9994 11468 11494
rect 11532 10674 11560 11698
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11150 11652 11562
rect 12256 11452 12552 11472
rect 12312 11450 12336 11452
rect 12392 11450 12416 11452
rect 12472 11450 12496 11452
rect 12334 11398 12336 11450
rect 12398 11398 12410 11450
rect 12472 11398 12474 11450
rect 12312 11396 12336 11398
rect 12392 11396 12416 11398
rect 12472 11396 12496 11398
rect 12256 11376 12552 11396
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10130 11560 10610
rect 11624 10470 11652 11086
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10520 9110 10548 9522
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9256 8188 9552 8208
rect 9312 8186 9336 8188
rect 9392 8186 9416 8188
rect 9472 8186 9496 8188
rect 9334 8134 9336 8186
rect 9398 8134 9410 8186
rect 9472 8134 9474 8186
rect 9312 8132 9336 8134
rect 9392 8132 9416 8134
rect 9472 8132 9496 8134
rect 9256 8112 9552 8132
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7886 8984 8026
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8680 7546 8708 7754
rect 8956 7546 8984 7822
rect 9876 7750 9904 8230
rect 9968 7954 9996 8434
rect 10060 8090 10088 8434
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 7756 6556 8052 6576
rect 7812 6554 7836 6556
rect 7892 6554 7916 6556
rect 7972 6554 7996 6556
rect 7834 6502 7836 6554
rect 7898 6502 7910 6554
rect 7972 6502 7974 6554
rect 7812 6500 7836 6502
rect 7892 6500 7916 6502
rect 7972 6500 7996 6502
rect 7756 6480 8052 6500
rect 8128 6118 8156 6734
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8588 5914 8616 6734
rect 8680 6322 8708 6734
rect 9140 6662 9168 7346
rect 9256 7100 9552 7120
rect 9312 7098 9336 7100
rect 9392 7098 9416 7100
rect 9472 7098 9496 7100
rect 9334 7046 9336 7098
rect 9398 7046 9410 7098
rect 9472 7046 9474 7098
rect 9312 7044 9336 7046
rect 9392 7044 9416 7046
rect 9472 7044 9496 7046
rect 9256 7024 9552 7044
rect 9876 6730 9904 7686
rect 9968 7342 9996 7890
rect 10060 7478 10088 8026
rect 10336 7750 10364 8910
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10336 7410 10364 7686
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 10520 6798 10548 9046
rect 10612 8498 10640 9522
rect 11440 9450 11468 9930
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11624 9382 11652 9930
rect 11716 9518 11744 10678
rect 11900 10470 11928 10950
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11900 9654 11928 10406
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 9178 11652 9318
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11900 8974 11928 9386
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 10756 8732 11052 8752
rect 10812 8730 10836 8732
rect 10892 8730 10916 8732
rect 10972 8730 10996 8732
rect 10834 8678 10836 8730
rect 10898 8678 10910 8730
rect 10972 8678 10974 8730
rect 10812 8676 10836 8678
rect 10892 8676 10916 8678
rect 10972 8676 10996 8678
rect 10756 8656 11052 8676
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11716 8090 11744 8434
rect 11900 8294 11928 8910
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 10756 7644 11052 7664
rect 10812 7642 10836 7644
rect 10892 7642 10916 7644
rect 10972 7642 10996 7644
rect 10834 7590 10836 7642
rect 10898 7590 10910 7642
rect 10972 7590 10974 7642
rect 10812 7588 10836 7590
rect 10892 7588 10916 7590
rect 10972 7588 10996 7590
rect 10756 7568 11052 7588
rect 11256 7546 11284 7686
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7656 5636 7708 5642
rect 7576 5596 7656 5624
rect 7656 5578 7708 5584
rect 7668 5370 7696 5578
rect 7756 5468 8052 5488
rect 7812 5466 7836 5468
rect 7892 5466 7916 5468
rect 7972 5466 7996 5468
rect 7834 5414 7836 5466
rect 7898 5414 7910 5466
rect 7972 5414 7974 5466
rect 7812 5412 7836 5414
rect 7892 5412 7916 5414
rect 7972 5412 7996 5414
rect 7756 5392 8052 5412
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 3256 4924 3552 4944
rect 3312 4922 3336 4924
rect 3392 4922 3416 4924
rect 3472 4922 3496 4924
rect 3334 4870 3336 4922
rect 3398 4870 3410 4922
rect 3472 4870 3474 4922
rect 3312 4868 3336 4870
rect 3392 4868 3416 4870
rect 3472 4868 3496 4870
rect 3256 4848 3552 4868
rect 6256 4924 6552 4944
rect 6312 4922 6336 4924
rect 6392 4922 6416 4924
rect 6472 4922 6496 4924
rect 6334 4870 6336 4922
rect 6398 4870 6410 4922
rect 6472 4870 6474 4922
rect 6312 4868 6336 4870
rect 6392 4868 6416 4870
rect 6472 4868 6496 4870
rect 6256 4848 6552 4868
rect 8128 4826 8156 5646
rect 8680 5370 8708 6258
rect 9140 6254 9168 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5710 9168 6190
rect 9256 6012 9552 6032
rect 9312 6010 9336 6012
rect 9392 6010 9416 6012
rect 9472 6010 9496 6012
rect 9334 5958 9336 6010
rect 9398 5958 9410 6010
rect 9472 5958 9474 6010
rect 9312 5956 9336 5958
rect 9392 5956 9416 5958
rect 9472 5956 9496 5958
rect 9256 5936 9552 5956
rect 9692 5846 9720 6394
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8852 5568 8904 5574
rect 8852 5510 8904 5516
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 1756 4380 2052 4400
rect 1812 4378 1836 4380
rect 1892 4378 1916 4380
rect 1972 4378 1996 4380
rect 1834 4326 1836 4378
rect 1898 4326 1910 4378
rect 1972 4326 1974 4378
rect 1812 4324 1836 4326
rect 1892 4324 1916 4326
rect 1972 4324 1996 4326
rect 1756 4304 2052 4324
rect 4756 4380 5052 4400
rect 4812 4378 4836 4380
rect 4892 4378 4916 4380
rect 4972 4378 4996 4380
rect 4834 4326 4836 4378
rect 4898 4326 4910 4378
rect 4972 4326 4974 4378
rect 4812 4324 4836 4326
rect 4892 4324 4916 4326
rect 4972 4324 4996 4326
rect 4756 4304 5052 4324
rect 7756 4380 8052 4400
rect 7812 4378 7836 4380
rect 7892 4378 7916 4380
rect 7972 4378 7996 4380
rect 7834 4326 7836 4378
rect 7898 4326 7910 4378
rect 7972 4326 7974 4378
rect 7812 4324 7836 4326
rect 7892 4324 7916 4326
rect 7972 4324 7996 4326
rect 7756 4304 8052 4324
rect 8220 4282 8248 4626
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8772 4146 8800 4966
rect 8864 4185 8892 5510
rect 9048 5370 9076 5578
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9692 5234 9720 5782
rect 9876 5642 9904 6666
rect 10520 6458 10548 6734
rect 11716 6662 11744 7346
rect 11900 6798 11928 8230
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 10756 6556 11052 6576
rect 10812 6554 10836 6556
rect 10892 6554 10916 6556
rect 10972 6554 10996 6556
rect 10834 6502 10836 6554
rect 10898 6502 10910 6554
rect 10972 6502 10974 6554
rect 10812 6500 10836 6502
rect 10892 6500 10916 6502
rect 10972 6500 10996 6502
rect 10756 6480 11052 6500
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 11164 6254 11192 6598
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 10520 5778 10548 6190
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 10060 5370 10088 5646
rect 11348 5642 11376 6326
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 10756 5468 11052 5488
rect 10812 5466 10836 5468
rect 10892 5466 10916 5468
rect 10972 5466 10996 5468
rect 10834 5414 10836 5466
rect 10898 5414 10910 5466
rect 10972 5414 10974 5466
rect 10812 5412 10836 5414
rect 10892 5412 10916 5414
rect 10972 5412 10996 5414
rect 10756 5392 11052 5412
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 8956 4486 8984 5170
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9256 4924 9552 4944
rect 9312 4922 9336 4924
rect 9392 4922 9416 4924
rect 9472 4922 9496 4924
rect 9334 4870 9336 4922
rect 9398 4870 9410 4922
rect 9472 4870 9474 4922
rect 9312 4868 9336 4870
rect 9392 4868 9416 4870
rect 9472 4868 9496 4870
rect 9256 4848 9552 4868
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8850 4176 8906 4185
rect 8116 4140 8168 4146
rect 8116 4082 8168 4088
rect 8760 4140 8812 4146
rect 8850 4111 8906 4120
rect 8760 4082 8812 4088
rect 3256 3836 3552 3856
rect 3312 3834 3336 3836
rect 3392 3834 3416 3836
rect 3472 3834 3496 3836
rect 3334 3782 3336 3834
rect 3398 3782 3410 3834
rect 3472 3782 3474 3834
rect 3312 3780 3336 3782
rect 3392 3780 3416 3782
rect 3472 3780 3496 3782
rect 3256 3760 3552 3780
rect 6256 3836 6552 3856
rect 6312 3834 6336 3836
rect 6392 3834 6416 3836
rect 6472 3834 6496 3836
rect 6334 3782 6336 3834
rect 6398 3782 6410 3834
rect 6472 3782 6474 3834
rect 6312 3780 6336 3782
rect 6392 3780 6416 3782
rect 6472 3780 6496 3782
rect 6256 3760 6552 3780
rect 8128 3670 8156 4082
rect 8668 4072 8720 4078
rect 8772 4049 8800 4082
rect 8864 4078 8892 4111
rect 8852 4072 8904 4078
rect 8668 4014 8720 4020
rect 8758 4040 8814 4049
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 1756 3292 2052 3312
rect 1812 3290 1836 3292
rect 1892 3290 1916 3292
rect 1972 3290 1996 3292
rect 1834 3238 1836 3290
rect 1898 3238 1910 3290
rect 1972 3238 1974 3290
rect 1812 3236 1836 3238
rect 1892 3236 1916 3238
rect 1972 3236 1996 3238
rect 1756 3216 2052 3236
rect 4756 3292 5052 3312
rect 4812 3290 4836 3292
rect 4892 3290 4916 3292
rect 4972 3290 4996 3292
rect 4834 3238 4836 3290
rect 4898 3238 4910 3290
rect 4972 3238 4974 3290
rect 4812 3236 4836 3238
rect 4892 3236 4916 3238
rect 4972 3236 4996 3238
rect 4756 3216 5052 3236
rect 7756 3292 8052 3312
rect 7812 3290 7836 3292
rect 7892 3290 7916 3292
rect 7972 3290 7996 3292
rect 7834 3238 7836 3290
rect 7898 3238 7910 3290
rect 7972 3238 7974 3290
rect 7812 3236 7836 3238
rect 7892 3236 7916 3238
rect 7972 3236 7996 3238
rect 7756 3216 8052 3236
rect 8680 3058 8708 4014
rect 8852 4014 8904 4020
rect 8758 3975 8814 3984
rect 8772 3738 8800 3975
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8772 3194 8800 3674
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 3256 2748 3552 2768
rect 3312 2746 3336 2748
rect 3392 2746 3416 2748
rect 3472 2746 3496 2748
rect 3334 2694 3336 2746
rect 3398 2694 3410 2746
rect 3472 2694 3474 2746
rect 3312 2692 3336 2694
rect 3392 2692 3416 2694
rect 3472 2692 3496 2694
rect 3256 2672 3552 2692
rect 6256 2748 6552 2768
rect 6312 2746 6336 2748
rect 6392 2746 6416 2748
rect 6472 2746 6496 2748
rect 6334 2694 6336 2746
rect 6398 2694 6410 2746
rect 6472 2694 6474 2746
rect 6312 2692 6336 2694
rect 6392 2692 6416 2694
rect 6472 2692 6496 2694
rect 6256 2672 6552 2692
rect 8680 2650 8708 2994
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8956 2446 8984 4422
rect 9692 4214 9720 4966
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9968 4126 10180 4154
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9772 4072 9824 4078
rect 9968 4049 9996 4126
rect 10152 4078 10180 4126
rect 10140 4072 10192 4078
rect 9772 4014 9824 4020
rect 9954 4040 10010 4049
rect 9140 3398 9168 4014
rect 9256 3836 9552 3856
rect 9312 3834 9336 3836
rect 9392 3834 9416 3836
rect 9472 3834 9496 3836
rect 9334 3782 9336 3834
rect 9398 3782 9410 3834
rect 9472 3782 9474 3834
rect 9312 3780 9336 3782
rect 9392 3780 9416 3782
rect 9472 3780 9496 3782
rect 9256 3760 9552 3780
rect 9784 3466 9812 4014
rect 10140 4014 10192 4020
rect 9954 3975 10010 3984
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 1756 2204 2052 2224
rect 1812 2202 1836 2204
rect 1892 2202 1916 2204
rect 1972 2202 1996 2204
rect 1834 2150 1836 2202
rect 1898 2150 1910 2202
rect 1972 2150 1974 2202
rect 1812 2148 1836 2150
rect 1892 2148 1916 2150
rect 1972 2148 1996 2150
rect 1756 2128 2052 2148
rect 4756 2204 5052 2224
rect 4812 2202 4836 2204
rect 4892 2202 4916 2204
rect 4972 2202 4996 2204
rect 4834 2150 4836 2202
rect 4898 2150 4910 2202
rect 4972 2150 4974 2202
rect 4812 2148 4836 2150
rect 4892 2148 4916 2150
rect 4972 2148 4996 2150
rect 4756 2128 5052 2148
rect 7756 2204 8052 2224
rect 7812 2202 7836 2204
rect 7892 2202 7916 2204
rect 7972 2202 7996 2204
rect 7834 2150 7836 2202
rect 7898 2150 7910 2202
rect 7972 2150 7974 2202
rect 7812 2148 7836 2150
rect 7892 2148 7916 2150
rect 7972 2148 7996 2150
rect 7756 2128 8052 2148
rect 296 1352 348 1358
rect 296 1294 348 1300
rect 18 82 74 800
rect 308 82 336 1294
rect 18 54 336 82
rect 9140 82 9168 3334
rect 9784 3126 9812 3402
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10152 3058 10180 4014
rect 10244 3738 10272 4558
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10244 3126 10272 3674
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 9256 2748 9552 2768
rect 9312 2746 9336 2748
rect 9392 2746 9416 2748
rect 9472 2746 9496 2748
rect 9334 2694 9336 2746
rect 9398 2694 9410 2746
rect 9472 2694 9474 2746
rect 9312 2692 9336 2694
rect 9392 2692 9416 2694
rect 9472 2692 9496 2694
rect 9256 2672 9552 2692
rect 10336 1358 10364 5306
rect 11348 5234 11376 5578
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11152 5228 11204 5234
rect 11336 5228 11388 5234
rect 11204 5188 11284 5216
rect 11152 5170 11204 5176
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11072 4826 11100 5102
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10416 4548 10468 4554
rect 10416 4490 10468 4496
rect 10428 3466 10456 4490
rect 10756 4380 11052 4400
rect 10812 4378 10836 4380
rect 10892 4378 10916 4380
rect 10972 4378 10996 4380
rect 10834 4326 10836 4378
rect 10898 4326 10910 4378
rect 10972 4326 10974 4378
rect 10812 4324 10836 4326
rect 10892 4324 10916 4326
rect 10972 4324 10996 4326
rect 10756 4304 11052 4324
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10428 2582 10456 3402
rect 10520 2854 10548 3402
rect 10756 3292 11052 3312
rect 10812 3290 10836 3292
rect 10892 3290 10916 3292
rect 10972 3290 10996 3292
rect 10834 3238 10836 3290
rect 10898 3238 10910 3290
rect 10972 3238 10974 3290
rect 10812 3236 10836 3238
rect 10892 3236 10916 3238
rect 10972 3236 10996 3238
rect 10756 3216 11052 3236
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10520 2650 10548 2790
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10796 2446 10824 2858
rect 10980 2446 11008 2926
rect 11164 2514 11192 5034
rect 11256 4214 11284 5188
rect 11336 5170 11388 5176
rect 11348 4758 11376 5170
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11440 4690 11468 5238
rect 11532 5166 11560 5646
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11716 5098 11744 6598
rect 11900 6118 11928 6734
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 5370 11836 5578
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11900 5250 11928 6054
rect 11992 5778 12020 10950
rect 12176 10810 12204 11086
rect 12636 11014 12664 11698
rect 12820 11354 12848 12038
rect 13280 11898 13308 12922
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13372 12646 13400 12718
rect 13464 12646 13492 13330
rect 13556 13190 13584 13806
rect 14016 13786 14136 13814
rect 14016 13394 14044 13786
rect 14384 13462 14412 13874
rect 15256 13628 15552 13648
rect 15312 13626 15336 13628
rect 15392 13626 15416 13628
rect 15472 13626 15496 13628
rect 15334 13574 15336 13626
rect 15398 13574 15410 13626
rect 15472 13574 15474 13626
rect 15312 13572 15336 13574
rect 15392 13572 15416 13574
rect 15472 13572 15496 13574
rect 15256 13552 15552 13572
rect 15580 13462 15608 13942
rect 15764 13938 15792 14962
rect 15948 14414 15976 15302
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15764 13530 15792 13874
rect 16132 13870 16160 15438
rect 16756 15260 17052 15280
rect 16812 15258 16836 15260
rect 16892 15258 16916 15260
rect 16972 15258 16996 15260
rect 16834 15206 16836 15258
rect 16898 15206 16910 15258
rect 16972 15206 16974 15258
rect 16812 15204 16836 15206
rect 16892 15204 16916 15206
rect 16972 15204 16996 15206
rect 16756 15184 17052 15204
rect 17420 14822 17448 15506
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17604 14890 17632 15438
rect 17696 14958 17724 15438
rect 17972 14958 18000 16186
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 18156 15502 18184 15982
rect 18256 15804 18552 15824
rect 18312 15802 18336 15804
rect 18392 15802 18416 15804
rect 18472 15802 18496 15804
rect 18334 15750 18336 15802
rect 18398 15750 18410 15802
rect 18472 15750 18474 15802
rect 18312 15748 18336 15750
rect 18392 15748 18416 15750
rect 18472 15748 18496 15750
rect 18256 15728 18552 15748
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 18156 15094 18184 15438
rect 19168 15094 19196 15438
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 19444 15026 19472 15506
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13556 11898 13584 13126
rect 13648 12442 13676 13330
rect 13756 13084 14052 13104
rect 13812 13082 13836 13084
rect 13892 13082 13916 13084
rect 13972 13082 13996 13084
rect 13834 13030 13836 13082
rect 13898 13030 13910 13082
rect 13972 13030 13974 13082
rect 13812 13028 13836 13030
rect 13892 13028 13916 13030
rect 13972 13028 13996 13030
rect 13756 13008 14052 13028
rect 14200 12850 14228 13330
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13188 11354 13216 11562
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13280 11218 13308 11834
rect 13648 11286 13676 12378
rect 13740 12170 13768 12718
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14292 12442 14320 12650
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13756 11996 14052 12016
rect 13812 11994 13836 11996
rect 13892 11994 13916 11996
rect 13972 11994 13996 11996
rect 13834 11942 13836 11994
rect 13898 11942 13910 11994
rect 13972 11942 13974 11994
rect 13812 11940 13836 11942
rect 13892 11940 13916 11942
rect 13972 11940 13996 11942
rect 13756 11920 14052 11940
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 13756 10908 14052 10928
rect 13812 10906 13836 10908
rect 13892 10906 13916 10908
rect 13972 10906 13996 10908
rect 13834 10854 13836 10906
rect 13898 10854 13910 10906
rect 13972 10854 13974 10906
rect 13812 10852 13836 10854
rect 13892 10852 13916 10854
rect 13972 10852 13996 10854
rect 13756 10832 14052 10852
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 14004 10600 14056 10606
rect 14108 10588 14136 11630
rect 14292 11286 14320 11766
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14292 11014 14320 11222
rect 14384 11218 14412 12582
rect 14568 11898 14596 13262
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 14844 12646 14872 13194
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14056 10560 14136 10588
rect 14004 10542 14056 10548
rect 12256 10364 12552 10384
rect 12312 10362 12336 10364
rect 12392 10362 12416 10364
rect 12472 10362 12496 10364
rect 12334 10310 12336 10362
rect 12398 10310 12410 10362
rect 12472 10310 12474 10362
rect 12312 10308 12336 10310
rect 12392 10308 12416 10310
rect 12472 10308 12496 10310
rect 12256 10288 12552 10308
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12256 9276 12552 9296
rect 12312 9274 12336 9276
rect 12392 9274 12416 9276
rect 12472 9274 12496 9276
rect 12334 9222 12336 9274
rect 12398 9222 12410 9274
rect 12472 9222 12474 9274
rect 12312 9220 12336 9222
rect 12392 9220 12416 9222
rect 12472 9220 12496 9222
rect 12256 9200 12552 9220
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 12728 8498 12756 8842
rect 12912 8838 12940 9522
rect 13556 9450 13584 10542
rect 14016 10266 14044 10542
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9722 13676 9998
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 13756 9820 14052 9840
rect 13812 9818 13836 9820
rect 13892 9818 13916 9820
rect 13972 9818 13996 9820
rect 13834 9766 13836 9818
rect 13898 9766 13910 9818
rect 13972 9766 13974 9818
rect 13812 9764 13836 9766
rect 13892 9764 13916 9766
rect 13972 9764 13996 9766
rect 13756 9744 14052 9764
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8566 12940 8774
rect 13756 8732 14052 8752
rect 13812 8730 13836 8732
rect 13892 8730 13916 8732
rect 13972 8730 13996 8732
rect 13834 8678 13836 8730
rect 13898 8678 13910 8730
rect 13972 8678 13974 8730
rect 13812 8676 13836 8678
rect 13892 8676 13916 8678
rect 13972 8676 13996 8678
rect 13756 8656 14052 8676
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12256 8188 12552 8208
rect 12312 8186 12336 8188
rect 12392 8186 12416 8188
rect 12472 8186 12496 8188
rect 12334 8134 12336 8186
rect 12398 8134 12410 8186
rect 12472 8134 12474 8186
rect 12312 8132 12336 8134
rect 12392 8132 12416 8134
rect 12472 8132 12496 8134
rect 12256 8112 12552 8132
rect 12728 8090 12756 8434
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12912 8022 12940 8502
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12912 7410 12940 7958
rect 13280 7954 13308 8366
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 14016 7886 14044 8230
rect 13820 7880 13872 7886
rect 13648 7840 13820 7868
rect 13648 7546 13676 7840
rect 13820 7822 13872 7828
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13756 7644 14052 7664
rect 13812 7642 13836 7644
rect 13892 7642 13916 7644
rect 13972 7642 13996 7644
rect 13834 7590 13836 7642
rect 13898 7590 13910 7642
rect 13972 7590 13974 7642
rect 13812 7588 13836 7590
rect 13892 7588 13916 7590
rect 13972 7588 13996 7590
rect 13756 7568 14052 7588
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11808 5222 11928 5250
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4214 11652 4558
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11612 4208 11664 4214
rect 11808 4185 11836 5222
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11612 4150 11664 4156
rect 11794 4176 11850 4185
rect 11256 4078 11284 4150
rect 11900 4146 11928 4490
rect 11992 4486 12020 5714
rect 12084 5234 12112 7142
rect 12256 7100 12552 7120
rect 12312 7098 12336 7100
rect 12392 7098 12416 7100
rect 12472 7098 12496 7100
rect 12334 7046 12336 7098
rect 12398 7046 12410 7098
rect 12472 7046 12474 7098
rect 12312 7044 12336 7046
rect 12392 7044 12416 7046
rect 12472 7044 12496 7046
rect 12256 7024 12552 7044
rect 12636 6866 12664 7278
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12636 6254 12664 6666
rect 12912 6390 12940 7142
rect 13096 6730 13124 7142
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13096 6458 13124 6666
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12256 6012 12552 6032
rect 12312 6010 12336 6012
rect 12392 6010 12416 6012
rect 12472 6010 12496 6012
rect 12334 5958 12336 6010
rect 12398 5958 12410 6010
rect 12472 5958 12474 6010
rect 12312 5956 12336 5958
rect 12392 5956 12416 5958
rect 12472 5956 12496 5958
rect 12256 5936 12552 5956
rect 12636 5914 12664 6190
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13004 5710 13032 6054
rect 13096 5914 13124 6258
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13096 5778 13124 5850
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13188 5710 13216 6802
rect 13464 6322 13492 7210
rect 13740 7002 13768 7346
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13756 6556 14052 6576
rect 13812 6554 13836 6556
rect 13892 6554 13916 6556
rect 13972 6554 13996 6556
rect 13834 6502 13836 6554
rect 13898 6502 13910 6554
rect 13972 6502 13974 6554
rect 13812 6500 13836 6502
rect 13892 6500 13916 6502
rect 13972 6500 13996 6502
rect 13756 6480 14052 6500
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12072 5228 12124 5234
rect 12124 5188 12204 5216
rect 12072 5170 12124 5176
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 12070 4176 12126 4185
rect 11794 4111 11850 4120
rect 11888 4140 11940 4146
rect 12070 4111 12126 4120
rect 11888 4082 11940 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 11256 2446 11284 3878
rect 11900 3738 11928 4082
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 12084 3194 12112 4111
rect 12176 3466 12204 5188
rect 13004 5166 13032 5646
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12256 4924 12552 4944
rect 12312 4922 12336 4924
rect 12392 4922 12416 4924
rect 12472 4922 12496 4924
rect 12334 4870 12336 4922
rect 12398 4870 12410 4922
rect 12472 4870 12474 4922
rect 12312 4868 12336 4870
rect 12392 4868 12416 4870
rect 12472 4868 12496 4870
rect 12256 4848 12552 4868
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12256 3836 12552 3856
rect 12312 3834 12336 3836
rect 12392 3834 12416 3836
rect 12472 3834 12496 3836
rect 12334 3782 12336 3834
rect 12398 3782 12410 3834
rect 12472 3782 12474 3834
rect 12312 3780 12336 3782
rect 12392 3780 12416 3782
rect 12472 3780 12496 3782
rect 12256 3760 12552 3780
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11348 2514 11376 2994
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 12084 2446 12112 3130
rect 12176 2514 12204 3402
rect 12636 3058 12664 4218
rect 13188 3942 13216 5646
rect 13756 5468 14052 5488
rect 13812 5466 13836 5468
rect 13892 5466 13916 5468
rect 13972 5466 13996 5468
rect 13834 5414 13836 5466
rect 13898 5414 13910 5466
rect 13972 5414 13974 5466
rect 13812 5412 13836 5414
rect 13892 5412 13916 5414
rect 13972 5412 13996 5414
rect 13756 5392 14052 5412
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13756 4380 14052 4400
rect 13812 4378 13836 4380
rect 13892 4378 13916 4380
rect 13972 4378 13996 4380
rect 13834 4326 13836 4378
rect 13898 4326 13910 4378
rect 13972 4326 13974 4378
rect 13812 4324 13836 4326
rect 13892 4324 13916 4326
rect 13972 4324 13996 4326
rect 13756 4304 14052 4324
rect 14108 4282 14136 9658
rect 14200 9450 14228 9862
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14292 9178 14320 10950
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14476 10198 14504 10678
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14568 9722 14596 11834
rect 14844 11286 14872 12582
rect 15120 12102 15148 13194
rect 15580 12986 15608 13398
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15856 12646 15884 13670
rect 16132 13394 16160 13806
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15256 12540 15552 12560
rect 15312 12538 15336 12540
rect 15392 12538 15416 12540
rect 15472 12538 15496 12540
rect 15334 12486 15336 12538
rect 15398 12486 15410 12538
rect 15472 12486 15474 12538
rect 15312 12484 15336 12486
rect 15392 12484 15416 12486
rect 15472 12484 15496 12486
rect 15256 12464 15552 12484
rect 15856 12306 15884 12582
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 11762 15148 12038
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14936 11354 14964 11698
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 15120 11082 15148 11698
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15256 11452 15552 11472
rect 15312 11450 15336 11452
rect 15392 11450 15416 11452
rect 15472 11450 15496 11452
rect 15334 11398 15336 11450
rect 15398 11398 15410 11450
rect 15472 11398 15474 11450
rect 15312 11396 15336 11398
rect 15392 11396 15416 11398
rect 15472 11396 15496 11398
rect 15256 11376 15552 11396
rect 15672 11150 15700 11630
rect 15948 11150 15976 12310
rect 16224 12238 16252 12718
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16224 11286 16252 12174
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15672 10674 15700 11086
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15256 10364 15552 10384
rect 15312 10362 15336 10364
rect 15392 10362 15416 10364
rect 15472 10362 15496 10364
rect 15334 10310 15336 10362
rect 15398 10310 15410 10362
rect 15472 10310 15474 10362
rect 15312 10308 15336 10310
rect 15392 10308 15416 10310
rect 15472 10308 15496 10310
rect 15256 10288 15552 10308
rect 15948 10266 15976 11086
rect 16040 10810 16068 11154
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 15672 9654 15700 10066
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14476 9178 14504 9522
rect 15256 9276 15552 9296
rect 15312 9274 15336 9276
rect 15392 9274 15416 9276
rect 15472 9274 15496 9276
rect 15334 9222 15336 9274
rect 15398 9222 15410 9274
rect 15472 9222 15474 9274
rect 15312 9220 15336 9222
rect 15392 9220 15416 9222
rect 15472 9220 15496 9222
rect 15256 9200 15552 9220
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7546 14320 7822
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14292 7274 14320 7482
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14200 5370 14228 6938
rect 14292 6866 14320 7210
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14384 6440 14412 8910
rect 14476 8430 14504 9114
rect 16040 9042 16068 10746
rect 16224 9722 16252 11222
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 8566 14964 8774
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14936 8090 14964 8502
rect 15120 8498 15148 8910
rect 15580 8634 15608 8910
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 8294 15148 8434
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 15120 7954 15148 8230
rect 15256 8188 15552 8208
rect 15312 8186 15336 8188
rect 15392 8186 15416 8188
rect 15472 8186 15496 8188
rect 15334 8134 15336 8186
rect 15398 8134 15410 8186
rect 15472 8134 15474 8186
rect 15312 8132 15336 8134
rect 15392 8132 15416 8134
rect 15472 8132 15496 8134
rect 15256 8112 15552 8132
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15580 7410 15608 8570
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15256 7100 15552 7120
rect 15312 7098 15336 7100
rect 15392 7098 15416 7100
rect 15472 7098 15496 7100
rect 15334 7046 15336 7098
rect 15398 7046 15410 7098
rect 15472 7046 15474 7098
rect 15312 7044 15336 7046
rect 15392 7044 15416 7046
rect 15472 7044 15496 7046
rect 15256 7024 15552 7044
rect 15580 6934 15608 7346
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 14384 6412 14504 6440
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14292 5574 14320 6190
rect 14384 6118 14412 6258
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 3126 13216 3334
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12256 2748 12552 2768
rect 12312 2746 12336 2748
rect 12392 2746 12416 2748
rect 12472 2746 12496 2748
rect 12334 2694 12336 2746
rect 12398 2694 12410 2746
rect 12472 2694 12474 2746
rect 12312 2692 12336 2694
rect 12392 2692 12416 2694
rect 12472 2692 12496 2694
rect 12256 2672 12552 2692
rect 13188 2650 13216 3062
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13556 2582 13584 4150
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13648 3738 13676 3878
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13648 3534 13676 3674
rect 14108 3602 14136 4014
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13756 3292 14052 3312
rect 13812 3290 13836 3292
rect 13892 3290 13916 3292
rect 13972 3290 13996 3292
rect 13834 3238 13836 3290
rect 13898 3238 13910 3290
rect 13972 3238 13974 3290
rect 13812 3236 13836 3238
rect 13892 3236 13916 3238
rect 13972 3236 13996 3238
rect 13756 3216 14052 3236
rect 14108 2990 14136 3538
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 13740 2854 13768 2926
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 13740 2446 13768 2790
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 11256 2310 11284 2382
rect 14200 2310 14228 4558
rect 14292 2650 14320 5510
rect 14384 5234 14412 6054
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 4486 14412 5170
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14384 2378 14412 4422
rect 14476 4214 14504 6412
rect 15256 6012 15552 6032
rect 15312 6010 15336 6012
rect 15392 6010 15416 6012
rect 15472 6010 15496 6012
rect 15334 5958 15336 6010
rect 15398 5958 15410 6010
rect 15472 5958 15474 6010
rect 15312 5956 15336 5958
rect 15392 5956 15416 5958
rect 15472 5956 15496 5958
rect 15256 5936 15552 5956
rect 15764 5914 15792 7686
rect 15856 7478 15884 7822
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 15856 6934 15884 7414
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15948 6730 15976 7142
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 6186 15976 6666
rect 16040 6322 16068 8842
rect 16132 7868 16160 9454
rect 16224 9178 16252 9658
rect 16316 9586 16344 11494
rect 16408 11218 16436 14282
rect 16684 13870 16712 14350
rect 16756 14172 17052 14192
rect 16812 14170 16836 14172
rect 16892 14170 16916 14172
rect 16972 14170 16996 14172
rect 16834 14118 16836 14170
rect 16898 14118 16910 14170
rect 16972 14118 16974 14170
rect 16812 14116 16836 14118
rect 16892 14116 16916 14118
rect 16972 14116 16996 14118
rect 16756 14096 17052 14116
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11762 16528 12174
rect 16592 11898 16620 12786
rect 16684 12782 16712 13806
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16756 13084 17052 13104
rect 16812 13082 16836 13084
rect 16892 13082 16916 13084
rect 16972 13082 16996 13084
rect 16834 13030 16836 13082
rect 16898 13030 16910 13082
rect 16972 13030 16974 13082
rect 16812 13028 16836 13030
rect 16892 13028 16916 13030
rect 16972 13028 16996 13030
rect 16756 13008 17052 13028
rect 17144 12986 17172 13262
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16684 12442 16712 12718
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16776 12322 16804 12786
rect 17132 12640 17184 12646
rect 17236 12628 17264 13330
rect 17184 12600 17264 12628
rect 17132 12582 17184 12588
rect 16684 12294 16804 12322
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16500 11354 16528 11698
rect 16684 11558 16712 12294
rect 16756 11996 17052 12016
rect 16812 11994 16836 11996
rect 16892 11994 16916 11996
rect 16972 11994 16996 11996
rect 16834 11942 16836 11994
rect 16898 11942 16910 11994
rect 16972 11942 16974 11994
rect 16812 11940 16836 11942
rect 16892 11940 16916 11942
rect 16972 11940 16996 11942
rect 16756 11920 17052 11940
rect 17144 11898 17172 12582
rect 17328 12238 17356 14010
rect 17420 13870 17448 14758
rect 17604 14618 17632 14826
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 14006 17632 14350
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17420 12850 17448 13806
rect 17604 13258 17632 13942
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17696 12442 17724 14894
rect 17972 14618 18000 14894
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18256 14716 18552 14736
rect 18312 14714 18336 14716
rect 18392 14714 18416 14716
rect 18472 14714 18496 14716
rect 18334 14662 18336 14714
rect 18398 14662 18410 14714
rect 18472 14662 18474 14714
rect 18312 14660 18336 14662
rect 18392 14660 18416 14662
rect 18472 14660 18496 14662
rect 18256 14640 18552 14660
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 12442 17816 14214
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 11898 17356 12174
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 10198 16436 11154
rect 16500 11150 16528 11290
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16500 10742 16528 11086
rect 17144 11014 17172 11698
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 16756 10908 17052 10928
rect 16812 10906 16836 10908
rect 16892 10906 16916 10908
rect 16972 10906 16996 10908
rect 16834 10854 16836 10906
rect 16898 10854 16910 10906
rect 16972 10854 16974 10906
rect 16812 10852 16836 10854
rect 16892 10852 16916 10854
rect 16972 10852 16996 10854
rect 16756 10832 17052 10852
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16776 10062 16804 10406
rect 16580 10056 16632 10062
rect 16764 10056 16816 10062
rect 16632 10016 16712 10044
rect 16580 9998 16632 10004
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16316 8498 16344 9386
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16304 8492 16356 8498
rect 16356 8452 16436 8480
rect 16304 8434 16356 8440
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 7880 16264 7886
rect 16132 7840 16212 7868
rect 16132 7546 16160 7840
rect 16212 7822 16264 7828
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16316 6866 16344 8230
rect 16408 7478 16436 8452
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14568 4826 14596 5646
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15120 5234 15148 5578
rect 15948 5556 15976 6122
rect 16040 5846 16068 6258
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 16028 5568 16080 5574
rect 15948 5528 16028 5556
rect 16028 5510 16080 5516
rect 16040 5302 16068 5510
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 15120 4690 15148 5170
rect 15256 4924 15552 4944
rect 15312 4922 15336 4924
rect 15392 4922 15416 4924
rect 15472 4922 15496 4924
rect 15334 4870 15336 4922
rect 15398 4870 15410 4922
rect 15472 4870 15474 4922
rect 15312 4868 15336 4870
rect 15392 4868 15416 4870
rect 15472 4868 15496 4870
rect 15256 4848 15552 4868
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 15396 4154 15424 4694
rect 16132 4690 16160 6054
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15396 4146 15608 4154
rect 15384 4140 15608 4146
rect 15436 4126 15608 4140
rect 15384 4082 15436 4088
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 15028 3398 15056 3878
rect 15256 3836 15552 3856
rect 15312 3834 15336 3836
rect 15392 3834 15416 3836
rect 15472 3834 15496 3836
rect 15334 3782 15336 3834
rect 15398 3782 15410 3834
rect 15472 3782 15474 3834
rect 15312 3780 15336 3782
rect 15392 3780 15416 3782
rect 15472 3780 15496 3782
rect 15256 3760 15552 3780
rect 15580 3670 15608 4126
rect 15856 3942 15884 4558
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 16132 3738 16160 4626
rect 16224 3942 16252 5510
rect 16316 5166 16344 6802
rect 16500 6662 16528 8978
rect 16592 8838 16620 9522
rect 16684 9382 16712 10016
rect 16764 9998 16816 10004
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 16756 9820 17052 9840
rect 16812 9818 16836 9820
rect 16892 9818 16916 9820
rect 16972 9818 16996 9820
rect 16834 9766 16836 9818
rect 16898 9766 16910 9818
rect 16972 9766 16974 9818
rect 16812 9764 16836 9766
rect 16892 9764 16916 9766
rect 16972 9764 16996 9766
rect 16756 9744 17052 9764
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 6866 16620 8774
rect 16684 7886 16712 9318
rect 17144 8974 17172 9862
rect 17328 9518 17356 9998
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17420 9042 17448 9862
rect 17604 9722 17632 10610
rect 17972 10470 18000 14554
rect 18892 13938 18920 14758
rect 18984 14414 19012 14826
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 18984 14074 19012 14350
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18256 13628 18552 13648
rect 18312 13626 18336 13628
rect 18392 13626 18416 13628
rect 18472 13626 18496 13628
rect 18334 13574 18336 13626
rect 18398 13574 18410 13626
rect 18472 13574 18474 13626
rect 18312 13572 18336 13574
rect 18392 13572 18416 13574
rect 18472 13572 18496 13574
rect 18256 13552 18552 13572
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18156 11898 18184 12718
rect 18256 12540 18552 12560
rect 18312 12538 18336 12540
rect 18392 12538 18416 12540
rect 18472 12538 18496 12540
rect 18334 12486 18336 12538
rect 18398 12486 18410 12538
rect 18472 12486 18474 12538
rect 18312 12484 18336 12486
rect 18392 12484 18416 12486
rect 18472 12484 18496 12486
rect 18256 12464 18552 12484
rect 18616 12374 18644 12854
rect 18708 12374 18736 13670
rect 18892 13530 18920 13874
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18604 11688 18656 11694
rect 18708 11676 18736 12310
rect 18800 12170 18828 13194
rect 19076 12986 19104 14214
rect 19444 14074 19472 14350
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19168 13462 19196 14010
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13462 19472 13806
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19536 13326 19564 15302
rect 19628 14414 19656 15982
rect 19904 15570 19932 16050
rect 21256 15804 21552 15824
rect 21312 15802 21336 15804
rect 21392 15802 21416 15804
rect 21472 15802 21496 15804
rect 21334 15750 21336 15802
rect 21398 15750 21410 15802
rect 21472 15750 21474 15802
rect 21312 15748 21336 15750
rect 21392 15748 21416 15750
rect 21472 15748 21496 15750
rect 21256 15728 21552 15748
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 19756 15260 20052 15280
rect 19812 15258 19836 15260
rect 19892 15258 19916 15260
rect 19972 15258 19996 15260
rect 19834 15206 19836 15258
rect 19898 15206 19910 15258
rect 19972 15206 19974 15258
rect 19812 15204 19836 15206
rect 19892 15204 19916 15206
rect 19972 15204 19996 15206
rect 19756 15184 20052 15204
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20180 14618 20208 14962
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19628 13870 19656 14214
rect 19756 14172 20052 14192
rect 19812 14170 19836 14172
rect 19892 14170 19916 14172
rect 19972 14170 19996 14172
rect 19834 14118 19836 14170
rect 19898 14118 19910 14170
rect 19972 14118 19974 14170
rect 19812 14116 19836 14118
rect 19892 14116 19916 14118
rect 19972 14116 19996 14118
rect 19756 14096 20052 14116
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 20076 13796 20128 13802
rect 20076 13738 20128 13744
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19536 12986 19564 13262
rect 19756 13084 20052 13104
rect 19812 13082 19836 13084
rect 19892 13082 19916 13084
rect 19972 13082 19996 13084
rect 19834 13030 19836 13082
rect 19898 13030 19910 13082
rect 19972 13030 19974 13082
rect 19812 13028 19836 13030
rect 19892 13028 19916 13030
rect 19972 13028 19996 13030
rect 19756 13008 20052 13028
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11898 18828 12106
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18656 11648 18736 11676
rect 18604 11630 18656 11636
rect 18256 11452 18552 11472
rect 18312 11450 18336 11452
rect 18392 11450 18416 11452
rect 18472 11450 18496 11452
rect 18334 11398 18336 11450
rect 18398 11398 18410 11450
rect 18472 11398 18474 11450
rect 18312 11396 18336 11398
rect 18392 11396 18416 11398
rect 18472 11396 18496 11398
rect 18256 11376 18552 11396
rect 18616 11014 18644 11630
rect 18892 11540 18920 12174
rect 19756 11996 20052 12016
rect 19812 11994 19836 11996
rect 19892 11994 19916 11996
rect 19972 11994 19996 11996
rect 19834 11942 19836 11994
rect 19898 11942 19910 11994
rect 19972 11942 19974 11994
rect 19812 11940 19836 11942
rect 19892 11940 19916 11942
rect 19972 11940 19996 11942
rect 19756 11920 20052 11940
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 18800 11512 18920 11540
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 18256 10364 18552 10384
rect 18312 10362 18336 10364
rect 18392 10362 18416 10364
rect 18472 10362 18496 10364
rect 18334 10310 18336 10362
rect 18398 10310 18410 10362
rect 18472 10310 18474 10362
rect 18312 10308 18336 10310
rect 18392 10308 18416 10310
rect 18472 10308 18496 10310
rect 18256 10288 18552 10308
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18248 9722 18276 9930
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18256 9276 18552 9296
rect 18312 9274 18336 9276
rect 18392 9274 18416 9276
rect 18472 9274 18496 9276
rect 18334 9222 18336 9274
rect 18398 9222 18410 9274
rect 18472 9222 18474 9274
rect 18312 9220 18336 9222
rect 18392 9220 18416 9222
rect 18472 9220 18496 9222
rect 18256 9200 18552 9220
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16756 8732 17052 8752
rect 16812 8730 16836 8732
rect 16892 8730 16916 8732
rect 16972 8730 16996 8732
rect 16834 8678 16836 8730
rect 16898 8678 16910 8730
rect 16972 8678 16974 8730
rect 16812 8676 16836 8678
rect 16892 8676 16916 8678
rect 16972 8676 16996 8678
rect 16756 8656 17052 8676
rect 17144 8634 17172 8910
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17420 8090 17448 8978
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 7206 16712 7822
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 17224 7812 17276 7818
rect 17224 7754 17276 7760
rect 16756 7644 17052 7664
rect 16812 7642 16836 7644
rect 16892 7642 16916 7644
rect 16972 7642 16996 7644
rect 16834 7590 16836 7642
rect 16898 7590 16910 7642
rect 16972 7590 16974 7642
rect 16812 7588 16836 7590
rect 16892 7588 16916 7590
rect 16972 7588 16996 7590
rect 16756 7568 17052 7588
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 17052 7002 17080 7346
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6322 16528 6598
rect 16756 6556 17052 6576
rect 16812 6554 16836 6556
rect 16892 6554 16916 6556
rect 16972 6554 16996 6556
rect 16834 6502 16836 6554
rect 16898 6502 16910 6554
rect 16972 6502 16974 6554
rect 16812 6500 16836 6502
rect 16892 6500 16916 6502
rect 16972 6500 16996 6502
rect 16756 6480 17052 6500
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16408 5030 16436 6190
rect 16500 5370 16528 6258
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 5370 16712 5646
rect 16756 5468 17052 5488
rect 16812 5466 16836 5468
rect 16892 5466 16916 5468
rect 16972 5466 16996 5468
rect 16834 5414 16836 5466
rect 16898 5414 16910 5466
rect 16972 5414 16974 5466
rect 16812 5412 16836 5414
rect 16892 5412 16916 5414
rect 16972 5412 16996 5414
rect 16756 5392 17052 5412
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4554 16436 4966
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16684 4214 16712 5306
rect 16756 4380 17052 4400
rect 16812 4378 16836 4380
rect 16892 4378 16916 4380
rect 16972 4378 16996 4380
rect 16834 4326 16836 4378
rect 16898 4326 16910 4378
rect 16972 4326 16974 4378
rect 16812 4324 16836 4326
rect 16892 4324 16916 4326
rect 16972 4324 16996 4326
rect 16756 4304 17052 4324
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14476 2650 14504 3062
rect 15028 2990 15056 3334
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 15028 2514 15056 2926
rect 15580 2922 15608 3606
rect 16224 3534 16252 3878
rect 17144 3584 17172 7754
rect 17236 7546 17264 7754
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17512 7410 17540 8230
rect 17880 7750 17908 8842
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18156 8090 18184 8434
rect 18256 8188 18552 8208
rect 18312 8186 18336 8188
rect 18392 8186 18416 8188
rect 18472 8186 18496 8188
rect 18334 8134 18336 8186
rect 18398 8134 18410 8186
rect 18472 8134 18474 8186
rect 18312 8132 18336 8134
rect 18392 8132 18416 8134
rect 18472 8132 18496 8134
rect 18256 8112 18552 8132
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18156 7886 18184 8026
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 18156 7546 18184 7822
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 18256 7100 18552 7120
rect 18312 7098 18336 7100
rect 18392 7098 18416 7100
rect 18472 7098 18496 7100
rect 18334 7046 18336 7098
rect 18398 7046 18410 7098
rect 18472 7046 18474 7098
rect 18312 7044 18336 7046
rect 18392 7044 18416 7046
rect 18472 7044 18496 7046
rect 18256 7024 18552 7044
rect 18616 6798 18644 10950
rect 18800 9926 18828 11512
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17604 6458 17632 6666
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17420 5710 17448 6326
rect 18156 6118 18184 6734
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5302 17632 5646
rect 18156 5302 18184 6054
rect 18256 6012 18552 6032
rect 18312 6010 18336 6012
rect 18392 6010 18416 6012
rect 18472 6010 18496 6012
rect 18334 5958 18336 6010
rect 18398 5958 18410 6010
rect 18472 5958 18474 6010
rect 18312 5956 18336 5958
rect 18392 5956 18416 5958
rect 18472 5956 18496 5958
rect 18256 5936 18552 5956
rect 18616 5574 18644 6190
rect 18708 5778 18736 7686
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17236 4010 17264 4558
rect 17420 4282 17448 5170
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17880 4690 17908 5102
rect 18156 4826 18184 5238
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18256 4924 18552 4944
rect 18312 4922 18336 4924
rect 18392 4922 18416 4924
rect 18472 4922 18496 4924
rect 18334 4870 18336 4922
rect 18398 4870 18410 4922
rect 18472 4870 18474 4922
rect 18312 4868 18336 4870
rect 18392 4868 18416 4870
rect 18472 4868 18496 4870
rect 18256 4848 18552 4868
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 18616 4622 18644 5170
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 18156 4146 18184 4558
rect 18708 4146 18736 5102
rect 18800 4554 18828 9862
rect 18984 9654 19012 10066
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 18984 8022 19012 9590
rect 19076 9382 19104 9998
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 8294 19104 9318
rect 19168 9042 19196 10610
rect 19260 10538 19288 11086
rect 19444 11082 19472 11698
rect 19720 11354 19748 11698
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11354 20024 11494
rect 19708 11348 19760 11354
rect 19628 11308 19708 11336
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19444 10810 19472 11018
rect 19628 10810 19656 11308
rect 19708 11290 19760 11296
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19756 10908 20052 10928
rect 19812 10906 19836 10908
rect 19892 10906 19916 10908
rect 19972 10906 19996 10908
rect 19834 10854 19836 10906
rect 19898 10854 19910 10906
rect 19972 10854 19974 10906
rect 19812 10852 19836 10854
rect 19892 10852 19916 10854
rect 19972 10852 19996 10854
rect 19756 10832 20052 10852
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19260 9994 19288 10474
rect 20088 10266 20116 13738
rect 20180 13734 20208 14350
rect 20272 14006 20300 14418
rect 20364 14074 20392 15030
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20272 13530 20300 13942
rect 20548 13870 20576 14282
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20548 13530 20576 13806
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20272 12782 20300 13466
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20180 12102 20208 12582
rect 20272 12442 20300 12718
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9586 19380 9862
rect 19340 9580 19392 9586
rect 19392 9540 19472 9568
rect 19340 9522 19392 9528
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19168 8498 19196 8978
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 8090 19104 8230
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18984 7002 19012 7958
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19076 6934 19104 8026
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19168 6866 19196 7346
rect 19156 6860 19208 6866
rect 19444 6848 19472 9540
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19536 8090 19564 9454
rect 19628 9178 19656 10066
rect 19756 9820 20052 9840
rect 19812 9818 19836 9820
rect 19892 9818 19916 9820
rect 19972 9818 19996 9820
rect 19834 9766 19836 9818
rect 19898 9766 19910 9818
rect 19972 9766 19974 9818
rect 19812 9764 19836 9766
rect 19892 9764 19916 9766
rect 19972 9764 19996 9766
rect 19756 9744 20052 9764
rect 20088 9586 20116 10202
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19720 9178 19748 9522
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19628 8498 19656 9114
rect 20180 8820 20208 12038
rect 20272 11762 20300 12378
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 10674 20484 11698
rect 20640 11558 20668 12786
rect 20732 11830 20760 15506
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 15162 21128 15438
rect 21272 15428 21324 15434
rect 21192 15388 21272 15416
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21100 14482 21128 15098
rect 21192 14958 21220 15388
rect 21272 15370 21324 15376
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21928 15162 21956 15370
rect 22756 15260 23052 15280
rect 22812 15258 22836 15260
rect 22892 15258 22916 15260
rect 22972 15258 22996 15260
rect 22834 15206 22836 15258
rect 22898 15206 22910 15258
rect 22972 15206 22974 15258
rect 22812 15204 22836 15206
rect 22892 15204 22916 15206
rect 22972 15204 22996 15206
rect 22756 15184 23052 15204
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21192 14618 21220 14894
rect 21256 14716 21552 14736
rect 21312 14714 21336 14716
rect 21392 14714 21416 14716
rect 21472 14714 21496 14716
rect 21334 14662 21336 14714
rect 21398 14662 21410 14714
rect 21472 14662 21474 14714
rect 21312 14660 21336 14662
rect 21392 14660 21416 14662
rect 21472 14660 21496 14662
rect 21256 14640 21552 14660
rect 21652 14618 21680 14962
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21652 14521 21680 14554
rect 21638 14512 21694 14521
rect 21088 14476 21140 14482
rect 21638 14447 21694 14456
rect 21916 14476 21968 14482
rect 21088 14418 21140 14424
rect 21916 14418 21968 14424
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21008 13530 21036 13874
rect 21928 13814 21956 14418
rect 23124 14346 23152 27338
rect 23216 27130 23244 27406
rect 25756 27228 26052 27248
rect 25812 27226 25836 27228
rect 25892 27226 25916 27228
rect 25972 27226 25996 27228
rect 25834 27174 25836 27226
rect 25898 27174 25910 27226
rect 25972 27174 25974 27226
rect 25812 27172 25836 27174
rect 25892 27172 25916 27174
rect 25972 27172 25996 27174
rect 25756 27152 26052 27172
rect 23204 27124 23256 27130
rect 23204 27066 23256 27072
rect 24256 26684 24552 26704
rect 24312 26682 24336 26684
rect 24392 26682 24416 26684
rect 24472 26682 24496 26684
rect 24334 26630 24336 26682
rect 24398 26630 24410 26682
rect 24472 26630 24474 26682
rect 24312 26628 24336 26630
rect 24392 26628 24416 26630
rect 24472 26628 24496 26630
rect 24256 26608 24552 26628
rect 27256 26684 27552 26704
rect 27312 26682 27336 26684
rect 27392 26682 27416 26684
rect 27472 26682 27496 26684
rect 27334 26630 27336 26682
rect 27398 26630 27410 26682
rect 27472 26630 27474 26682
rect 27312 26628 27336 26630
rect 27392 26628 27416 26630
rect 27472 26628 27496 26630
rect 27256 26608 27552 26628
rect 25756 26140 26052 26160
rect 25812 26138 25836 26140
rect 25892 26138 25916 26140
rect 25972 26138 25996 26140
rect 25834 26086 25836 26138
rect 25898 26086 25910 26138
rect 25972 26086 25974 26138
rect 25812 26084 25836 26086
rect 25892 26084 25916 26086
rect 25972 26084 25996 26086
rect 25756 26064 26052 26084
rect 24256 25596 24552 25616
rect 24312 25594 24336 25596
rect 24392 25594 24416 25596
rect 24472 25594 24496 25596
rect 24334 25542 24336 25594
rect 24398 25542 24410 25594
rect 24472 25542 24474 25594
rect 24312 25540 24336 25542
rect 24392 25540 24416 25542
rect 24472 25540 24496 25542
rect 24256 25520 24552 25540
rect 27256 25596 27552 25616
rect 27312 25594 27336 25596
rect 27392 25594 27416 25596
rect 27472 25594 27496 25596
rect 27334 25542 27336 25594
rect 27398 25542 27410 25594
rect 27472 25542 27474 25594
rect 27312 25540 27336 25542
rect 27392 25540 27416 25542
rect 27472 25540 27496 25542
rect 27256 25520 27552 25540
rect 25756 25052 26052 25072
rect 25812 25050 25836 25052
rect 25892 25050 25916 25052
rect 25972 25050 25996 25052
rect 25834 24998 25836 25050
rect 25898 24998 25910 25050
rect 25972 24998 25974 25050
rect 25812 24996 25836 24998
rect 25892 24996 25916 24998
rect 25972 24996 25996 24998
rect 25756 24976 26052 24996
rect 24256 24508 24552 24528
rect 24312 24506 24336 24508
rect 24392 24506 24416 24508
rect 24472 24506 24496 24508
rect 24334 24454 24336 24506
rect 24398 24454 24410 24506
rect 24472 24454 24474 24506
rect 24312 24452 24336 24454
rect 24392 24452 24416 24454
rect 24472 24452 24496 24454
rect 24256 24432 24552 24452
rect 27256 24508 27552 24528
rect 27312 24506 27336 24508
rect 27392 24506 27416 24508
rect 27472 24506 27496 24508
rect 27334 24454 27336 24506
rect 27398 24454 27410 24506
rect 27472 24454 27474 24506
rect 27312 24452 27336 24454
rect 27392 24452 27416 24454
rect 27472 24452 27496 24454
rect 27256 24432 27552 24452
rect 25756 23964 26052 23984
rect 25812 23962 25836 23964
rect 25892 23962 25916 23964
rect 25972 23962 25996 23964
rect 25834 23910 25836 23962
rect 25898 23910 25910 23962
rect 25972 23910 25974 23962
rect 25812 23908 25836 23910
rect 25892 23908 25916 23910
rect 25972 23908 25996 23910
rect 25756 23888 26052 23908
rect 24256 23420 24552 23440
rect 24312 23418 24336 23420
rect 24392 23418 24416 23420
rect 24472 23418 24496 23420
rect 24334 23366 24336 23418
rect 24398 23366 24410 23418
rect 24472 23366 24474 23418
rect 24312 23364 24336 23366
rect 24392 23364 24416 23366
rect 24472 23364 24496 23366
rect 24256 23344 24552 23364
rect 27256 23420 27552 23440
rect 27312 23418 27336 23420
rect 27392 23418 27416 23420
rect 27472 23418 27496 23420
rect 27334 23366 27336 23418
rect 27398 23366 27410 23418
rect 27472 23366 27474 23418
rect 27312 23364 27336 23366
rect 27392 23364 27416 23366
rect 27472 23364 27496 23366
rect 27256 23344 27552 23364
rect 25756 22876 26052 22896
rect 25812 22874 25836 22876
rect 25892 22874 25916 22876
rect 25972 22874 25996 22876
rect 25834 22822 25836 22874
rect 25898 22822 25910 22874
rect 25972 22822 25974 22874
rect 25812 22820 25836 22822
rect 25892 22820 25916 22822
rect 25972 22820 25996 22822
rect 25756 22800 26052 22820
rect 24256 22332 24552 22352
rect 24312 22330 24336 22332
rect 24392 22330 24416 22332
rect 24472 22330 24496 22332
rect 24334 22278 24336 22330
rect 24398 22278 24410 22330
rect 24472 22278 24474 22330
rect 24312 22276 24336 22278
rect 24392 22276 24416 22278
rect 24472 22276 24496 22278
rect 24256 22256 24552 22276
rect 27256 22332 27552 22352
rect 27312 22330 27336 22332
rect 27392 22330 27416 22332
rect 27472 22330 27496 22332
rect 27334 22278 27336 22330
rect 27398 22278 27410 22330
rect 27472 22278 27474 22330
rect 27312 22276 27336 22278
rect 27392 22276 27416 22278
rect 27472 22276 27496 22278
rect 27256 22256 27552 22276
rect 25756 21788 26052 21808
rect 25812 21786 25836 21788
rect 25892 21786 25916 21788
rect 25972 21786 25996 21788
rect 25834 21734 25836 21786
rect 25898 21734 25910 21786
rect 25972 21734 25974 21786
rect 25812 21732 25836 21734
rect 25892 21732 25916 21734
rect 25972 21732 25996 21734
rect 25756 21712 26052 21732
rect 24256 21244 24552 21264
rect 24312 21242 24336 21244
rect 24392 21242 24416 21244
rect 24472 21242 24496 21244
rect 24334 21190 24336 21242
rect 24398 21190 24410 21242
rect 24472 21190 24474 21242
rect 24312 21188 24336 21190
rect 24392 21188 24416 21190
rect 24472 21188 24496 21190
rect 24256 21168 24552 21188
rect 27256 21244 27552 21264
rect 27312 21242 27336 21244
rect 27392 21242 27416 21244
rect 27472 21242 27496 21244
rect 27334 21190 27336 21242
rect 27398 21190 27410 21242
rect 27472 21190 27474 21242
rect 27312 21188 27336 21190
rect 27392 21188 27416 21190
rect 27472 21188 27496 21190
rect 27256 21168 27552 21188
rect 25756 20700 26052 20720
rect 25812 20698 25836 20700
rect 25892 20698 25916 20700
rect 25972 20698 25996 20700
rect 25834 20646 25836 20698
rect 25898 20646 25910 20698
rect 25972 20646 25974 20698
rect 25812 20644 25836 20646
rect 25892 20644 25916 20646
rect 25972 20644 25996 20646
rect 25756 20624 26052 20644
rect 24256 20156 24552 20176
rect 24312 20154 24336 20156
rect 24392 20154 24416 20156
rect 24472 20154 24496 20156
rect 24334 20102 24336 20154
rect 24398 20102 24410 20154
rect 24472 20102 24474 20154
rect 24312 20100 24336 20102
rect 24392 20100 24416 20102
rect 24472 20100 24496 20102
rect 24256 20080 24552 20100
rect 27256 20156 27552 20176
rect 27312 20154 27336 20156
rect 27392 20154 27416 20156
rect 27472 20154 27496 20156
rect 27334 20102 27336 20154
rect 27398 20102 27410 20154
rect 27472 20102 27474 20154
rect 27312 20100 27336 20102
rect 27392 20100 27416 20102
rect 27472 20100 27496 20102
rect 27256 20080 27552 20100
rect 25756 19612 26052 19632
rect 25812 19610 25836 19612
rect 25892 19610 25916 19612
rect 25972 19610 25996 19612
rect 25834 19558 25836 19610
rect 25898 19558 25910 19610
rect 25972 19558 25974 19610
rect 25812 19556 25836 19558
rect 25892 19556 25916 19558
rect 25972 19556 25996 19558
rect 25756 19536 26052 19556
rect 24256 19068 24552 19088
rect 24312 19066 24336 19068
rect 24392 19066 24416 19068
rect 24472 19066 24496 19068
rect 24334 19014 24336 19066
rect 24398 19014 24410 19066
rect 24472 19014 24474 19066
rect 24312 19012 24336 19014
rect 24392 19012 24416 19014
rect 24472 19012 24496 19014
rect 24256 18992 24552 19012
rect 27256 19068 27552 19088
rect 27312 19066 27336 19068
rect 27392 19066 27416 19068
rect 27472 19066 27496 19068
rect 27334 19014 27336 19066
rect 27398 19014 27410 19066
rect 27472 19014 27474 19066
rect 27312 19012 27336 19014
rect 27392 19012 27416 19014
rect 27472 19012 27496 19014
rect 27256 18992 27552 19012
rect 25756 18524 26052 18544
rect 25812 18522 25836 18524
rect 25892 18522 25916 18524
rect 25972 18522 25996 18524
rect 25834 18470 25836 18522
rect 25898 18470 25910 18522
rect 25972 18470 25974 18522
rect 25812 18468 25836 18470
rect 25892 18468 25916 18470
rect 25972 18468 25996 18470
rect 25756 18448 26052 18468
rect 24256 17980 24552 18000
rect 24312 17978 24336 17980
rect 24392 17978 24416 17980
rect 24472 17978 24496 17980
rect 24334 17926 24336 17978
rect 24398 17926 24410 17978
rect 24472 17926 24474 17978
rect 24312 17924 24336 17926
rect 24392 17924 24416 17926
rect 24472 17924 24496 17926
rect 24256 17904 24552 17924
rect 27256 17980 27552 18000
rect 27312 17978 27336 17980
rect 27392 17978 27416 17980
rect 27472 17978 27496 17980
rect 27334 17926 27336 17978
rect 27398 17926 27410 17978
rect 27472 17926 27474 17978
rect 27312 17924 27336 17926
rect 27392 17924 27416 17926
rect 27472 17924 27496 17926
rect 27256 17904 27552 17924
rect 25756 17436 26052 17456
rect 25812 17434 25836 17436
rect 25892 17434 25916 17436
rect 25972 17434 25996 17436
rect 25834 17382 25836 17434
rect 25898 17382 25910 17434
rect 25972 17382 25974 17434
rect 25812 17380 25836 17382
rect 25892 17380 25916 17382
rect 25972 17380 25996 17382
rect 25756 17360 26052 17380
rect 24256 16892 24552 16912
rect 24312 16890 24336 16892
rect 24392 16890 24416 16892
rect 24472 16890 24496 16892
rect 24334 16838 24336 16890
rect 24398 16838 24410 16890
rect 24472 16838 24474 16890
rect 24312 16836 24336 16838
rect 24392 16836 24416 16838
rect 24472 16836 24496 16838
rect 24256 16816 24552 16836
rect 27256 16892 27552 16912
rect 27312 16890 27336 16892
rect 27392 16890 27416 16892
rect 27472 16890 27496 16892
rect 27334 16838 27336 16890
rect 27398 16838 27410 16890
rect 27472 16838 27474 16890
rect 27312 16836 27336 16838
rect 27392 16836 27416 16838
rect 27472 16836 27496 16838
rect 27256 16816 27552 16836
rect 25756 16348 26052 16368
rect 25812 16346 25836 16348
rect 25892 16346 25916 16348
rect 25972 16346 25996 16348
rect 25834 16294 25836 16346
rect 25898 16294 25910 16346
rect 25972 16294 25974 16346
rect 25812 16292 25836 16294
rect 25892 16292 25916 16294
rect 25972 16292 25996 16294
rect 25756 16272 26052 16292
rect 24256 15804 24552 15824
rect 24312 15802 24336 15804
rect 24392 15802 24416 15804
rect 24472 15802 24496 15804
rect 24334 15750 24336 15802
rect 24398 15750 24410 15802
rect 24472 15750 24474 15802
rect 24312 15748 24336 15750
rect 24392 15748 24416 15750
rect 24472 15748 24496 15750
rect 24256 15728 24552 15748
rect 27256 15804 27552 15824
rect 27312 15802 27336 15804
rect 27392 15802 27416 15804
rect 27472 15802 27496 15804
rect 27334 15750 27336 15802
rect 27398 15750 27410 15802
rect 27472 15750 27474 15802
rect 27312 15748 27336 15750
rect 27392 15748 27416 15750
rect 27472 15748 27496 15750
rect 27256 15728 27552 15748
rect 25756 15260 26052 15280
rect 25812 15258 25836 15260
rect 25892 15258 25916 15260
rect 25972 15258 25996 15260
rect 25834 15206 25836 15258
rect 25898 15206 25910 15258
rect 25972 15206 25974 15258
rect 25812 15204 25836 15206
rect 25892 15204 25916 15206
rect 25972 15204 25996 15206
rect 25756 15184 26052 15204
rect 24256 14716 24552 14736
rect 24312 14714 24336 14716
rect 24392 14714 24416 14716
rect 24472 14714 24496 14716
rect 24334 14662 24336 14714
rect 24398 14662 24410 14714
rect 24472 14662 24474 14714
rect 24312 14660 24336 14662
rect 24392 14660 24416 14662
rect 24472 14660 24496 14662
rect 24256 14640 24552 14660
rect 27256 14716 27552 14736
rect 27312 14714 27336 14716
rect 27392 14714 27416 14716
rect 27472 14714 27496 14716
rect 27334 14662 27336 14714
rect 27398 14662 27410 14714
rect 27472 14662 27474 14714
rect 27312 14660 27336 14662
rect 27392 14660 27416 14662
rect 27472 14660 27496 14662
rect 27256 14640 27552 14660
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 21928 13802 22140 13814
rect 21928 13796 22152 13802
rect 21928 13786 22100 13796
rect 21256 13628 21552 13648
rect 21312 13626 21336 13628
rect 21392 13626 21416 13628
rect 21472 13626 21496 13628
rect 21334 13574 21336 13626
rect 21398 13574 21410 13626
rect 21472 13574 21474 13626
rect 21312 13572 21336 13574
rect 21392 13572 21416 13574
rect 21472 13572 21496 13574
rect 21256 13552 21552 13572
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21008 11830 21036 13126
rect 21100 12646 21128 13262
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21256 12540 21552 12560
rect 21312 12538 21336 12540
rect 21392 12538 21416 12540
rect 21472 12538 21496 12540
rect 21334 12486 21336 12538
rect 21398 12486 21410 12538
rect 21472 12486 21474 12538
rect 21312 12484 21336 12486
rect 21392 12484 21416 12486
rect 21472 12484 21496 12486
rect 21256 12464 21552 12484
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21100 11830 21128 12174
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20732 10810 20760 11766
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20364 10266 20392 10542
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20824 9654 20852 10610
rect 21008 10266 21036 11766
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 21100 11014 21128 11630
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21256 11452 21552 11472
rect 21312 11450 21336 11452
rect 21392 11450 21416 11452
rect 21472 11450 21496 11452
rect 21334 11398 21336 11450
rect 21398 11398 21410 11450
rect 21472 11398 21474 11450
rect 21312 11396 21336 11398
rect 21392 11396 21416 11398
rect 21472 11396 21496 11398
rect 21256 11376 21552 11396
rect 21836 11286 21864 11494
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21088 11008 21140 11014
rect 21088 10950 21140 10956
rect 21100 10742 21128 10950
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21192 10266 21220 10474
rect 21652 10470 21680 11086
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21256 10364 21552 10384
rect 21312 10362 21336 10364
rect 21392 10362 21416 10364
rect 21472 10362 21496 10364
rect 21334 10310 21336 10362
rect 21398 10310 21410 10362
rect 21472 10310 21474 10362
rect 21312 10308 21336 10310
rect 21392 10308 21416 10310
rect 21472 10308 21496 10310
rect 21256 10288 21552 10308
rect 20996 10260 21048 10266
rect 21180 10260 21232 10266
rect 20996 10202 21048 10208
rect 21100 10220 21180 10248
rect 20994 10024 21050 10033
rect 20994 9959 21050 9968
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20260 8832 20312 8838
rect 20180 8792 20260 8820
rect 20260 8774 20312 8780
rect 19756 8732 20052 8752
rect 19812 8730 19836 8732
rect 19892 8730 19916 8732
rect 19972 8730 19996 8732
rect 19834 8678 19836 8730
rect 19898 8678 19910 8730
rect 19972 8678 19974 8730
rect 19812 8676 19836 8678
rect 19892 8676 19916 8678
rect 19972 8676 19996 8678
rect 19756 8656 20052 8676
rect 20272 8498 20300 8774
rect 20824 8566 20852 9590
rect 21008 9586 21036 9959
rect 21100 9586 21128 10220
rect 21180 10202 21232 10208
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21100 9042 21128 9522
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 21192 8974 21220 9386
rect 21256 9276 21552 9296
rect 21312 9274 21336 9276
rect 21392 9274 21416 9276
rect 21472 9274 21496 9276
rect 21334 9222 21336 9274
rect 21398 9222 21410 9274
rect 21472 9222 21474 9274
rect 21312 9220 21336 9222
rect 21392 9220 21416 9222
rect 21472 9220 21496 9222
rect 21256 9200 21552 9220
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21192 8634 21220 8910
rect 21652 8650 21680 10406
rect 21928 10062 21956 13786
rect 22100 13738 22152 13744
rect 22664 13734 22692 14282
rect 22756 14172 23052 14192
rect 22812 14170 22836 14172
rect 22892 14170 22916 14172
rect 22972 14170 22996 14172
rect 22834 14118 22836 14170
rect 22898 14118 22910 14170
rect 22972 14118 22974 14170
rect 22812 14116 22836 14118
rect 22892 14116 22916 14118
rect 22972 14116 22996 14118
rect 22756 14096 23052 14116
rect 23124 14074 23152 14282
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23860 13814 23888 14418
rect 25756 14172 26052 14192
rect 25812 14170 25836 14172
rect 25892 14170 25916 14172
rect 25972 14170 25996 14172
rect 25834 14118 25836 14170
rect 25898 14118 25910 14170
rect 25972 14118 25974 14170
rect 25812 14116 25836 14118
rect 25892 14116 25916 14118
rect 25972 14116 25996 14118
rect 25756 14096 26052 14116
rect 23768 13786 23888 13814
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22020 12102 22048 12786
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22388 12238 22416 12718
rect 22572 12238 22600 12786
rect 22664 12374 22692 13670
rect 23768 13190 23796 13786
rect 24256 13628 24552 13648
rect 24312 13626 24336 13628
rect 24392 13626 24416 13628
rect 24472 13626 24496 13628
rect 24334 13574 24336 13626
rect 24398 13574 24410 13626
rect 24472 13574 24474 13626
rect 24312 13572 24336 13574
rect 24392 13572 24416 13574
rect 24472 13572 24496 13574
rect 24256 13552 24552 13572
rect 27256 13628 27552 13648
rect 27312 13626 27336 13628
rect 27392 13626 27416 13628
rect 27472 13626 27496 13628
rect 27334 13574 27336 13626
rect 27398 13574 27410 13626
rect 27472 13574 27474 13626
rect 27312 13572 27336 13574
rect 27392 13572 27416 13574
rect 27472 13572 27496 13574
rect 27256 13552 27552 13572
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 22756 13084 23052 13104
rect 22812 13082 22836 13084
rect 22892 13082 22916 13084
rect 22972 13082 22996 13084
rect 22834 13030 22836 13082
rect 22898 13030 22910 13082
rect 22972 13030 22974 13082
rect 22812 13028 22836 13030
rect 22892 13028 22916 13030
rect 22972 13028 22996 13030
rect 22756 13008 23052 13028
rect 23202 12744 23258 12753
rect 23768 12714 23796 13126
rect 25756 13084 26052 13104
rect 25812 13082 25836 13084
rect 25892 13082 25916 13084
rect 25972 13082 25996 13084
rect 25834 13030 25836 13082
rect 25898 13030 25910 13082
rect 25972 13030 25974 13082
rect 25812 13028 25836 13030
rect 25892 13028 25916 13030
rect 25972 13028 25996 13030
rect 25756 13008 26052 13028
rect 23202 12679 23258 12688
rect 23756 12708 23808 12714
rect 23216 12646 23244 12679
rect 23756 12650 23808 12656
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 23216 12442 23244 12582
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 22652 12368 22704 12374
rect 22652 12310 22704 12316
rect 23768 12238 23796 12650
rect 24256 12540 24552 12560
rect 24312 12538 24336 12540
rect 24392 12538 24416 12540
rect 24472 12538 24496 12540
rect 24334 12486 24336 12538
rect 24398 12486 24410 12538
rect 24472 12486 24474 12538
rect 24312 12484 24336 12486
rect 24392 12484 24416 12486
rect 24472 12484 24496 12486
rect 24256 12464 24552 12484
rect 27256 12540 27552 12560
rect 27312 12538 27336 12540
rect 27392 12538 27416 12540
rect 27472 12538 27496 12540
rect 27334 12486 27336 12538
rect 27398 12486 27410 12538
rect 27472 12486 27474 12538
rect 27312 12484 27336 12486
rect 27392 12484 27416 12486
rect 27472 12484 27496 12486
rect 27256 12464 27552 12484
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 22020 11558 22048 12038
rect 22388 11898 22416 12174
rect 22376 11892 22428 11898
rect 22376 11834 22428 11840
rect 22572 11762 22600 12174
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22020 11354 22048 11494
rect 22664 11354 22692 12174
rect 22756 11996 23052 12016
rect 22812 11994 22836 11996
rect 22892 11994 22916 11996
rect 22972 11994 22996 11996
rect 22834 11942 22836 11994
rect 22898 11942 22910 11994
rect 22972 11942 22974 11994
rect 22812 11940 22836 11942
rect 22892 11940 22916 11942
rect 22972 11940 22996 11942
rect 22756 11920 23052 11940
rect 25756 11996 26052 12016
rect 25812 11994 25836 11996
rect 25892 11994 25916 11996
rect 25972 11994 25996 11996
rect 25834 11942 25836 11994
rect 25898 11942 25910 11994
rect 25972 11942 25974 11994
rect 25812 11940 25836 11942
rect 25892 11940 25916 11942
rect 25972 11940 25996 11942
rect 25756 11920 26052 11940
rect 24256 11452 24552 11472
rect 24312 11450 24336 11452
rect 24392 11450 24416 11452
rect 24472 11450 24496 11452
rect 24334 11398 24336 11450
rect 24398 11398 24410 11450
rect 24472 11398 24474 11450
rect 24312 11396 24336 11398
rect 24392 11396 24416 11398
rect 24472 11396 24496 11398
rect 24256 11376 24552 11396
rect 27256 11452 27552 11472
rect 27312 11450 27336 11452
rect 27392 11450 27416 11452
rect 27472 11450 27496 11452
rect 27334 11398 27336 11450
rect 27398 11398 27410 11450
rect 27472 11398 27474 11450
rect 27312 11396 27336 11398
rect 27392 11396 27416 11398
rect 27472 11396 27496 11398
rect 27256 11376 27552 11396
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22480 10810 22508 11154
rect 28736 11121 28764 12310
rect 28722 11112 28778 11121
rect 28722 11047 28778 11056
rect 22756 10908 23052 10928
rect 22812 10906 22836 10908
rect 22892 10906 22916 10908
rect 22972 10906 22996 10908
rect 22834 10854 22836 10906
rect 22898 10854 22910 10906
rect 22972 10854 22974 10906
rect 22812 10852 22836 10854
rect 22892 10852 22916 10854
rect 22972 10852 22996 10854
rect 22756 10832 23052 10852
rect 25756 10908 26052 10928
rect 25812 10906 25836 10908
rect 25892 10906 25916 10908
rect 25972 10906 25996 10908
rect 25834 10854 25836 10906
rect 25898 10854 25910 10906
rect 25972 10854 25974 10906
rect 25812 10852 25836 10854
rect 25892 10852 25916 10854
rect 25972 10852 25996 10854
rect 25756 10832 26052 10852
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21560 8622 21680 8650
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 19628 8090 19656 8434
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 19628 7954 19656 8026
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19628 7546 19656 7890
rect 19904 7818 19932 8434
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19756 7644 20052 7664
rect 19812 7642 19836 7644
rect 19892 7642 19916 7644
rect 19972 7642 19996 7644
rect 19834 7590 19836 7642
rect 19898 7590 19910 7642
rect 19972 7590 19974 7642
rect 19812 7588 19836 7590
rect 19892 7588 19916 7590
rect 19972 7588 19996 7590
rect 19756 7568 20052 7588
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 20088 6866 20116 8366
rect 20272 8022 20300 8434
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20272 7002 20300 7958
rect 20456 7750 20484 8434
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20548 6866 20576 7142
rect 19524 6860 19576 6866
rect 19444 6820 19524 6848
rect 19156 6802 19208 6808
rect 19524 6802 19576 6808
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18892 5778 18920 6598
rect 19076 6390 19104 6598
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19076 5914 19104 6326
rect 19168 6254 19196 6802
rect 19340 6792 19392 6798
rect 19260 6752 19340 6780
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18892 4826 18920 5714
rect 19168 5710 19196 6190
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19168 5166 19196 5646
rect 19260 5642 19288 6752
rect 19340 6734 19392 6740
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19260 5370 19288 5578
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 19536 4282 19564 6802
rect 19756 6556 20052 6576
rect 19812 6554 19836 6556
rect 19892 6554 19916 6556
rect 19972 6554 19996 6556
rect 19834 6502 19836 6554
rect 19898 6502 19910 6554
rect 19972 6502 19974 6554
rect 19812 6500 19836 6502
rect 19892 6500 19916 6502
rect 19972 6500 19996 6502
rect 19756 6480 20052 6500
rect 20088 6458 20116 6802
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19812 5914 19840 6326
rect 19800 5908 19852 5914
rect 19628 5868 19800 5896
rect 19628 4826 19656 5868
rect 19800 5850 19852 5856
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 19756 5468 20052 5488
rect 19812 5466 19836 5468
rect 19892 5466 19916 5468
rect 19972 5466 19996 5468
rect 19834 5414 19836 5466
rect 19898 5414 19910 5466
rect 19972 5414 19974 5466
rect 19812 5412 19836 5414
rect 19892 5412 19916 5414
rect 19972 5412 19996 5414
rect 19756 5392 20052 5412
rect 20272 5302 20300 5850
rect 20640 5370 20668 7278
rect 20916 5778 20944 7346
rect 21008 5914 21036 7346
rect 21192 7342 21220 8570
rect 21560 8498 21588 8622
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21256 8188 21552 8208
rect 21312 8186 21336 8188
rect 21392 8186 21416 8188
rect 21472 8186 21496 8188
rect 21334 8134 21336 8186
rect 21398 8134 21410 8186
rect 21472 8134 21474 8186
rect 21312 8132 21336 8134
rect 21392 8132 21416 8134
rect 21472 8132 21496 8134
rect 21256 8112 21552 8132
rect 21652 7954 21680 8502
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21100 5914 21128 6802
rect 21192 6798 21220 7142
rect 21256 7100 21552 7120
rect 21312 7098 21336 7100
rect 21392 7098 21416 7100
rect 21472 7098 21496 7100
rect 21334 7046 21336 7098
rect 21398 7046 21410 7098
rect 21472 7046 21474 7098
rect 21312 7044 21336 7046
rect 21392 7044 21416 7046
rect 21472 7044 21496 7046
rect 21256 7024 21552 7044
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21192 6118 21220 6734
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 6458 21588 6666
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21652 6390 21680 7890
rect 21744 7886 21772 9930
rect 21928 9382 21956 9998
rect 21916 9376 21968 9382
rect 21916 9318 21968 9324
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21836 8090 21864 8910
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21744 7546 21772 7822
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21836 7478 21864 7754
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21744 6848 21772 7346
rect 21928 7206 21956 9318
rect 22020 8974 22048 10474
rect 24256 10364 24552 10384
rect 24312 10362 24336 10364
rect 24392 10362 24416 10364
rect 24472 10362 24496 10364
rect 24334 10310 24336 10362
rect 24398 10310 24410 10362
rect 24472 10310 24474 10362
rect 24312 10308 24336 10310
rect 24392 10308 24416 10310
rect 24472 10308 24496 10310
rect 24256 10288 24552 10308
rect 27256 10364 27552 10384
rect 27312 10362 27336 10364
rect 27392 10362 27416 10364
rect 27472 10362 27496 10364
rect 27334 10310 27336 10362
rect 27398 10310 27410 10362
rect 27472 10310 27474 10362
rect 27312 10308 27336 10310
rect 27392 10308 27416 10310
rect 27472 10308 27496 10310
rect 27256 10288 27552 10308
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 22296 9722 22324 9930
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22664 9722 22692 9862
rect 22756 9820 23052 9840
rect 22812 9818 22836 9820
rect 22892 9818 22916 9820
rect 22972 9818 22996 9820
rect 22834 9766 22836 9818
rect 22898 9766 22910 9818
rect 22972 9766 22974 9818
rect 22812 9764 22836 9766
rect 22892 9764 22916 9766
rect 22972 9764 22996 9766
rect 22756 9744 23052 9764
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 22020 8634 22048 8910
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22204 7392 22232 9386
rect 22296 9178 22324 9658
rect 24044 9586 24072 9930
rect 25756 9820 26052 9840
rect 25812 9818 25836 9820
rect 25892 9818 25916 9820
rect 25972 9818 25996 9820
rect 25834 9766 25836 9818
rect 25898 9766 25910 9818
rect 25972 9766 25974 9818
rect 25812 9764 25836 9766
rect 25892 9764 25916 9766
rect 25972 9764 25996 9766
rect 25756 9744 26052 9764
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22664 8634 22692 9522
rect 24256 9276 24552 9296
rect 24312 9274 24336 9276
rect 24392 9274 24416 9276
rect 24472 9274 24496 9276
rect 24334 9222 24336 9274
rect 24398 9222 24410 9274
rect 24472 9222 24474 9274
rect 24312 9220 24336 9222
rect 24392 9220 24416 9222
rect 24472 9220 24496 9222
rect 24256 9200 24552 9220
rect 27256 9276 27552 9296
rect 27312 9274 27336 9276
rect 27392 9274 27416 9276
rect 27472 9274 27496 9276
rect 27334 9222 27336 9274
rect 27398 9222 27410 9274
rect 27472 9222 27474 9274
rect 27312 9220 27336 9222
rect 27392 9220 27416 9222
rect 27472 9220 27496 9222
rect 27256 9200 27552 9220
rect 22756 8732 23052 8752
rect 22812 8730 22836 8732
rect 22892 8730 22916 8732
rect 22972 8730 22996 8732
rect 22834 8678 22836 8730
rect 22898 8678 22910 8730
rect 22972 8678 22974 8730
rect 22812 8676 22836 8678
rect 22892 8676 22916 8678
rect 22972 8676 22996 8678
rect 22756 8656 23052 8676
rect 25756 8732 26052 8752
rect 25812 8730 25836 8732
rect 25892 8730 25916 8732
rect 25972 8730 25996 8732
rect 25834 8678 25836 8730
rect 25898 8678 25910 8730
rect 25972 8678 25974 8730
rect 25812 8676 25836 8678
rect 25892 8676 25916 8678
rect 25972 8676 25996 8678
rect 25756 8656 26052 8676
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22480 8090 22508 8230
rect 24256 8188 24552 8208
rect 24312 8186 24336 8188
rect 24392 8186 24416 8188
rect 24472 8186 24496 8188
rect 24334 8134 24336 8186
rect 24398 8134 24410 8186
rect 24472 8134 24474 8186
rect 24312 8132 24336 8134
rect 24392 8132 24416 8134
rect 24472 8132 24496 8134
rect 24256 8112 24552 8132
rect 27256 8188 27552 8208
rect 27312 8186 27336 8188
rect 27392 8186 27416 8188
rect 27472 8186 27496 8188
rect 27334 8134 27336 8186
rect 27398 8134 27410 8186
rect 27472 8134 27474 8186
rect 27312 8132 27336 8134
rect 27392 8132 27416 8134
rect 27472 8132 27496 8134
rect 27256 8112 27552 8132
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22756 7644 23052 7664
rect 22812 7642 22836 7644
rect 22892 7642 22916 7644
rect 22972 7642 22996 7644
rect 22834 7590 22836 7642
rect 22898 7590 22910 7642
rect 22972 7590 22974 7642
rect 22812 7588 22836 7590
rect 22892 7588 22916 7590
rect 22972 7588 22996 7590
rect 22756 7568 23052 7588
rect 25756 7644 26052 7664
rect 25812 7642 25836 7644
rect 25892 7642 25916 7644
rect 25972 7642 25996 7644
rect 25834 7590 25836 7642
rect 25898 7590 25910 7642
rect 25972 7590 25974 7642
rect 25812 7588 25836 7590
rect 25892 7588 25916 7590
rect 25972 7588 25996 7590
rect 25756 7568 26052 7588
rect 22284 7404 22336 7410
rect 22204 7364 22284 7392
rect 22284 7346 22336 7352
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21824 6860 21876 6866
rect 21744 6820 21824 6848
rect 21640 6384 21692 6390
rect 21640 6326 21692 6332
rect 21744 6322 21772 6820
rect 21824 6802 21876 6808
rect 22296 6458 22324 7346
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 6730 22508 7142
rect 24256 7100 24552 7120
rect 24312 7098 24336 7100
rect 24392 7098 24416 7100
rect 24472 7098 24496 7100
rect 24334 7046 24336 7098
rect 24398 7046 24410 7098
rect 24472 7046 24474 7098
rect 24312 7044 24336 7046
rect 24392 7044 24416 7046
rect 24472 7044 24496 7046
rect 24256 7024 24552 7044
rect 27256 7100 27552 7120
rect 27312 7098 27336 7100
rect 27392 7098 27416 7100
rect 27472 7098 27496 7100
rect 27334 7046 27336 7098
rect 27398 7046 27410 7098
rect 27472 7046 27474 7098
rect 27312 7044 27336 7046
rect 27392 7044 27416 7046
rect 27472 7044 27496 7046
rect 27256 7024 27552 7044
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21256 6012 21552 6032
rect 21312 6010 21336 6012
rect 21392 6010 21416 6012
rect 21472 6010 21496 6012
rect 21334 5958 21336 6010
rect 21398 5958 21410 6010
rect 21472 5958 21474 6010
rect 21312 5956 21336 5958
rect 21392 5956 21416 5958
rect 21472 5956 21496 5958
rect 21256 5936 21552 5956
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20916 5370 20944 5714
rect 21744 5370 21772 6258
rect 22480 5914 22508 6666
rect 22756 6556 23052 6576
rect 22812 6554 22836 6556
rect 22892 6554 22916 6556
rect 22972 6554 22996 6556
rect 22834 6502 22836 6554
rect 22898 6502 22910 6554
rect 22972 6502 22974 6554
rect 22812 6500 22836 6502
rect 22892 6500 22916 6502
rect 22972 6500 22996 6502
rect 22756 6480 23052 6500
rect 25756 6556 26052 6576
rect 25812 6554 25836 6556
rect 25892 6554 25916 6556
rect 25972 6554 25996 6556
rect 25834 6502 25836 6554
rect 25898 6502 25910 6554
rect 25972 6502 25974 6554
rect 25812 6500 25836 6502
rect 25892 6500 25916 6502
rect 25972 6500 25996 6502
rect 25756 6480 26052 6500
rect 24256 6012 24552 6032
rect 24312 6010 24336 6012
rect 24392 6010 24416 6012
rect 24472 6010 24496 6012
rect 24334 5958 24336 6010
rect 24398 5958 24410 6010
rect 24472 5958 24474 6010
rect 24312 5956 24336 5958
rect 24392 5956 24416 5958
rect 24472 5956 24496 5958
rect 24256 5936 24552 5956
rect 27256 6012 27552 6032
rect 27312 6010 27336 6012
rect 27392 6010 27416 6012
rect 27472 6010 27496 6012
rect 27334 5958 27336 6010
rect 27398 5958 27410 6010
rect 27472 5958 27474 6010
rect 27312 5956 27336 5958
rect 27392 5956 27416 5958
rect 27472 5956 27496 5958
rect 27256 5936 27552 5956
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20180 4826 20208 5170
rect 21928 5166 21956 5510
rect 22756 5468 23052 5488
rect 22812 5466 22836 5468
rect 22892 5466 22916 5468
rect 22972 5466 22996 5468
rect 22834 5414 22836 5466
rect 22898 5414 22910 5466
rect 22972 5414 22974 5466
rect 22812 5412 22836 5414
rect 22892 5412 22916 5414
rect 22972 5412 22996 5414
rect 22756 5392 23052 5412
rect 25756 5468 26052 5488
rect 25812 5466 25836 5468
rect 25892 5466 25916 5468
rect 25972 5466 25996 5468
rect 25834 5414 25836 5466
rect 25898 5414 25910 5466
rect 25972 5414 25974 5466
rect 25812 5412 25836 5414
rect 25892 5412 25916 5414
rect 25972 5412 25996 5414
rect 25756 5392 26052 5412
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19628 4146 19656 4558
rect 19756 4380 20052 4400
rect 19812 4378 19836 4380
rect 19892 4378 19916 4380
rect 19972 4378 19996 4380
rect 19834 4326 19836 4378
rect 19898 4326 19910 4378
rect 19972 4326 19974 4378
rect 19812 4324 19836 4326
rect 19892 4324 19916 4326
rect 19972 4324 19996 4326
rect 19756 4304 20052 4324
rect 20456 4282 20484 5102
rect 21256 4924 21552 4944
rect 21312 4922 21336 4924
rect 21392 4922 21416 4924
rect 21472 4922 21496 4924
rect 21334 4870 21336 4922
rect 21398 4870 21410 4922
rect 21472 4870 21474 4922
rect 21312 4868 21336 4870
rect 21392 4868 21416 4870
rect 21472 4868 21496 4870
rect 21256 4848 21552 4868
rect 24256 4924 24552 4944
rect 24312 4922 24336 4924
rect 24392 4922 24416 4924
rect 24472 4922 24496 4924
rect 24334 4870 24336 4922
rect 24398 4870 24410 4922
rect 24472 4870 24474 4922
rect 24312 4868 24336 4870
rect 24392 4868 24416 4870
rect 24472 4868 24496 4870
rect 24256 4848 24552 4868
rect 27256 4924 27552 4944
rect 27312 4922 27336 4924
rect 27392 4922 27416 4924
rect 27472 4922 27496 4924
rect 27334 4870 27336 4922
rect 27398 4870 27410 4922
rect 27472 4870 27474 4922
rect 27312 4868 27336 4870
rect 27392 4868 27416 4870
rect 27472 4868 27496 4870
rect 27256 4848 27552 4868
rect 22756 4380 23052 4400
rect 22812 4378 22836 4380
rect 22892 4378 22916 4380
rect 22972 4378 22996 4380
rect 22834 4326 22836 4378
rect 22898 4326 22910 4378
rect 22972 4326 22974 4378
rect 22812 4324 22836 4326
rect 22892 4324 22916 4326
rect 22972 4324 22996 4326
rect 22756 4304 23052 4324
rect 25756 4380 26052 4400
rect 25812 4378 25836 4380
rect 25892 4378 25916 4380
rect 25972 4378 25996 4380
rect 25834 4326 25836 4378
rect 25898 4326 25910 4378
rect 25972 4326 25974 4378
rect 25812 4324 25836 4326
rect 25892 4324 25916 4326
rect 25972 4324 25996 4326
rect 25756 4304 26052 4324
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 18156 3602 18184 4082
rect 18256 3836 18552 3856
rect 18312 3834 18336 3836
rect 18392 3834 18416 3836
rect 18472 3834 18496 3836
rect 18334 3782 18336 3834
rect 18398 3782 18410 3834
rect 18472 3782 18474 3834
rect 18312 3780 18336 3782
rect 18392 3780 18416 3782
rect 18472 3780 18496 3782
rect 18256 3760 18552 3780
rect 18708 3738 18736 4082
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 17224 3596 17276 3602
rect 17144 3556 17224 3584
rect 17224 3538 17276 3544
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 16224 2854 16252 3470
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16316 2854 16344 3402
rect 16756 3292 17052 3312
rect 16812 3290 16836 3292
rect 16892 3290 16916 3292
rect 16972 3290 16996 3292
rect 16834 3238 16836 3290
rect 16898 3238 16910 3290
rect 16972 3238 16974 3290
rect 16812 3236 16836 3238
rect 16892 3236 16916 3238
rect 16972 3236 16996 3238
rect 16756 3216 17052 3236
rect 17236 3194 17264 3538
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 15256 2748 15552 2768
rect 15312 2746 15336 2748
rect 15392 2746 15416 2748
rect 15472 2746 15496 2748
rect 15334 2694 15336 2746
rect 15398 2694 15410 2746
rect 15472 2694 15474 2746
rect 15312 2692 15336 2694
rect 15392 2692 15416 2694
rect 15472 2692 15496 2694
rect 15256 2672 15552 2692
rect 16684 2514 16712 2994
rect 17788 2650 17816 3402
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 18156 2378 18184 2994
rect 18616 2922 18644 3470
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18256 2748 18552 2768
rect 18312 2746 18336 2748
rect 18392 2746 18416 2748
rect 18472 2746 18496 2748
rect 18334 2694 18336 2746
rect 18398 2694 18410 2746
rect 18472 2694 18474 2746
rect 18312 2692 18336 2694
rect 18392 2692 18416 2694
rect 18472 2692 18496 2694
rect 18256 2672 18552 2692
rect 18616 2446 18644 2858
rect 18708 2514 18736 3674
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 3194 19104 3538
rect 19628 3534 19656 4082
rect 21256 3836 21552 3856
rect 21312 3834 21336 3836
rect 21392 3834 21416 3836
rect 21472 3834 21496 3836
rect 21334 3782 21336 3834
rect 21398 3782 21410 3834
rect 21472 3782 21474 3834
rect 21312 3780 21336 3782
rect 21392 3780 21416 3782
rect 21472 3780 21496 3782
rect 21256 3760 21552 3780
rect 24256 3836 24552 3856
rect 24312 3834 24336 3836
rect 24392 3834 24416 3836
rect 24472 3834 24496 3836
rect 24334 3782 24336 3834
rect 24398 3782 24410 3834
rect 24472 3782 24474 3834
rect 24312 3780 24336 3782
rect 24392 3780 24416 3782
rect 24472 3780 24496 3782
rect 24256 3760 24552 3780
rect 27256 3836 27552 3856
rect 27312 3834 27336 3836
rect 27392 3834 27416 3836
rect 27472 3834 27496 3836
rect 27334 3782 27336 3834
rect 27398 3782 27410 3834
rect 27472 3782 27474 3834
rect 27312 3780 27336 3782
rect 27392 3780 27416 3782
rect 27472 3780 27496 3782
rect 27256 3760 27552 3780
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19756 3292 20052 3312
rect 19812 3290 19836 3292
rect 19892 3290 19916 3292
rect 19972 3290 19996 3292
rect 19834 3238 19836 3290
rect 19898 3238 19910 3290
rect 19972 3238 19974 3290
rect 19812 3236 19836 3238
rect 19892 3236 19916 3238
rect 19972 3236 19996 3238
rect 19756 3216 20052 3236
rect 22756 3292 23052 3312
rect 22812 3290 22836 3292
rect 22892 3290 22916 3292
rect 22972 3290 22996 3292
rect 22834 3238 22836 3290
rect 22898 3238 22910 3290
rect 22972 3238 22974 3290
rect 22812 3236 22836 3238
rect 22892 3236 22916 3238
rect 22972 3236 22996 3238
rect 22756 3216 23052 3236
rect 25756 3292 26052 3312
rect 25812 3290 25836 3292
rect 25892 3290 25916 3292
rect 25972 3290 25996 3292
rect 25834 3238 25836 3290
rect 25898 3238 25910 3290
rect 25972 3238 25974 3290
rect 25812 3236 25836 3238
rect 25892 3236 25916 3238
rect 25972 3236 25996 3238
rect 25756 3216 26052 3236
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 21256 2748 21552 2768
rect 21312 2746 21336 2748
rect 21392 2746 21416 2748
rect 21472 2746 21496 2748
rect 21334 2694 21336 2746
rect 21398 2694 21410 2746
rect 21472 2694 21474 2746
rect 21312 2692 21336 2694
rect 21392 2692 21416 2694
rect 21472 2692 21496 2694
rect 21256 2672 21552 2692
rect 24256 2748 24552 2768
rect 24312 2746 24336 2748
rect 24392 2746 24416 2748
rect 24472 2746 24496 2748
rect 24334 2694 24336 2746
rect 24398 2694 24410 2746
rect 24472 2694 24474 2746
rect 24312 2692 24336 2694
rect 24392 2692 24416 2694
rect 24472 2692 24496 2694
rect 24256 2672 24552 2692
rect 27256 2748 27552 2768
rect 27312 2746 27336 2748
rect 27392 2746 27416 2748
rect 27472 2746 27496 2748
rect 27334 2694 27336 2746
rect 27398 2694 27410 2746
rect 27472 2694 27474 2746
rect 27312 2692 27336 2694
rect 27392 2692 27416 2694
rect 27472 2692 27496 2694
rect 27256 2672 27552 2692
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 18144 2372 18196 2378
rect 18144 2314 18196 2320
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 10756 2204 11052 2224
rect 10812 2202 10836 2204
rect 10892 2202 10916 2204
rect 10972 2202 10996 2204
rect 10834 2150 10836 2202
rect 10898 2150 10910 2202
rect 10972 2150 10974 2202
rect 10812 2148 10836 2150
rect 10892 2148 10916 2150
rect 10972 2148 10996 2150
rect 10756 2128 11052 2148
rect 13756 2204 14052 2224
rect 13812 2202 13836 2204
rect 13892 2202 13916 2204
rect 13972 2202 13996 2204
rect 13834 2150 13836 2202
rect 13898 2150 13910 2202
rect 13972 2150 13974 2202
rect 13812 2148 13836 2150
rect 13892 2148 13916 2150
rect 13972 2148 13996 2150
rect 13756 2128 14052 2148
rect 16756 2204 17052 2224
rect 16812 2202 16836 2204
rect 16892 2202 16916 2204
rect 16972 2202 16996 2204
rect 16834 2150 16836 2202
rect 16898 2150 16910 2202
rect 16972 2150 16974 2202
rect 16812 2148 16836 2150
rect 16892 2148 16916 2150
rect 16972 2148 16996 2150
rect 16756 2128 17052 2148
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 9218 82 9274 800
rect 9140 54 9274 82
rect 18248 82 18276 2382
rect 19756 2204 20052 2224
rect 19812 2202 19836 2204
rect 19892 2202 19916 2204
rect 19972 2202 19996 2204
rect 19834 2150 19836 2202
rect 19898 2150 19910 2202
rect 19972 2150 19974 2202
rect 19812 2148 19836 2150
rect 19892 2148 19916 2150
rect 19972 2148 19996 2150
rect 19756 2128 20052 2148
rect 22756 2204 23052 2224
rect 22812 2202 22836 2204
rect 22892 2202 22916 2204
rect 22972 2202 22996 2204
rect 22834 2150 22836 2202
rect 22898 2150 22910 2202
rect 22972 2150 22974 2202
rect 22812 2148 22836 2150
rect 22892 2148 22916 2150
rect 22972 2148 22996 2150
rect 22756 2128 23052 2148
rect 25756 2204 26052 2224
rect 25812 2202 25836 2204
rect 25892 2202 25916 2204
rect 25972 2202 25996 2204
rect 25834 2150 25836 2202
rect 25898 2150 25910 2202
rect 25972 2150 25974 2202
rect 25812 2148 25836 2150
rect 25892 2148 25916 2150
rect 25972 2148 25996 2150
rect 25756 2128 26052 2148
rect 18510 82 18566 800
rect 18248 54 18566 82
rect 18 0 74 54
rect 9218 0 9274 54
rect 18510 0 18566 54
rect 27710 0 27766 800
<< via2 >>
rect 1756 29402 1812 29404
rect 1836 29402 1892 29404
rect 1916 29402 1972 29404
rect 1996 29402 2052 29404
rect 1756 29350 1782 29402
rect 1782 29350 1812 29402
rect 1836 29350 1846 29402
rect 1846 29350 1892 29402
rect 1916 29350 1962 29402
rect 1962 29350 1972 29402
rect 1996 29350 2026 29402
rect 2026 29350 2052 29402
rect 1756 29348 1812 29350
rect 1836 29348 1892 29350
rect 1916 29348 1972 29350
rect 1996 29348 2052 29350
rect 4756 29402 4812 29404
rect 4836 29402 4892 29404
rect 4916 29402 4972 29404
rect 4996 29402 5052 29404
rect 4756 29350 4782 29402
rect 4782 29350 4812 29402
rect 4836 29350 4846 29402
rect 4846 29350 4892 29402
rect 4916 29350 4962 29402
rect 4962 29350 4972 29402
rect 4996 29350 5026 29402
rect 5026 29350 5052 29402
rect 4756 29348 4812 29350
rect 4836 29348 4892 29350
rect 4916 29348 4972 29350
rect 4996 29348 5052 29350
rect 7756 29402 7812 29404
rect 7836 29402 7892 29404
rect 7916 29402 7972 29404
rect 7996 29402 8052 29404
rect 7756 29350 7782 29402
rect 7782 29350 7812 29402
rect 7836 29350 7846 29402
rect 7846 29350 7892 29402
rect 7916 29350 7962 29402
rect 7962 29350 7972 29402
rect 7996 29350 8026 29402
rect 8026 29350 8052 29402
rect 7756 29348 7812 29350
rect 7836 29348 7892 29350
rect 7916 29348 7972 29350
rect 7996 29348 8052 29350
rect 10756 29402 10812 29404
rect 10836 29402 10892 29404
rect 10916 29402 10972 29404
rect 10996 29402 11052 29404
rect 10756 29350 10782 29402
rect 10782 29350 10812 29402
rect 10836 29350 10846 29402
rect 10846 29350 10892 29402
rect 10916 29350 10962 29402
rect 10962 29350 10972 29402
rect 10996 29350 11026 29402
rect 11026 29350 11052 29402
rect 10756 29348 10812 29350
rect 10836 29348 10892 29350
rect 10916 29348 10972 29350
rect 10996 29348 11052 29350
rect 13756 29402 13812 29404
rect 13836 29402 13892 29404
rect 13916 29402 13972 29404
rect 13996 29402 14052 29404
rect 13756 29350 13782 29402
rect 13782 29350 13812 29402
rect 13836 29350 13846 29402
rect 13846 29350 13892 29402
rect 13916 29350 13962 29402
rect 13962 29350 13972 29402
rect 13996 29350 14026 29402
rect 14026 29350 14052 29402
rect 13756 29348 13812 29350
rect 13836 29348 13892 29350
rect 13916 29348 13972 29350
rect 13996 29348 14052 29350
rect 16756 29402 16812 29404
rect 16836 29402 16892 29404
rect 16916 29402 16972 29404
rect 16996 29402 17052 29404
rect 16756 29350 16782 29402
rect 16782 29350 16812 29402
rect 16836 29350 16846 29402
rect 16846 29350 16892 29402
rect 16916 29350 16962 29402
rect 16962 29350 16972 29402
rect 16996 29350 17026 29402
rect 17026 29350 17052 29402
rect 16756 29348 16812 29350
rect 16836 29348 16892 29350
rect 16916 29348 16972 29350
rect 16996 29348 17052 29350
rect 19756 29402 19812 29404
rect 19836 29402 19892 29404
rect 19916 29402 19972 29404
rect 19996 29402 20052 29404
rect 19756 29350 19782 29402
rect 19782 29350 19812 29402
rect 19836 29350 19846 29402
rect 19846 29350 19892 29402
rect 19916 29350 19962 29402
rect 19962 29350 19972 29402
rect 19996 29350 20026 29402
rect 20026 29350 20052 29402
rect 19756 29348 19812 29350
rect 19836 29348 19892 29350
rect 19916 29348 19972 29350
rect 19996 29348 20052 29350
rect 22756 29402 22812 29404
rect 22836 29402 22892 29404
rect 22916 29402 22972 29404
rect 22996 29402 23052 29404
rect 22756 29350 22782 29402
rect 22782 29350 22812 29402
rect 22836 29350 22846 29402
rect 22846 29350 22892 29402
rect 22916 29350 22962 29402
rect 22962 29350 22972 29402
rect 22996 29350 23026 29402
rect 23026 29350 23052 29402
rect 22756 29348 22812 29350
rect 22836 29348 22892 29350
rect 22916 29348 22972 29350
rect 22996 29348 23052 29350
rect 3256 28858 3312 28860
rect 3336 28858 3392 28860
rect 3416 28858 3472 28860
rect 3496 28858 3552 28860
rect 3256 28806 3282 28858
rect 3282 28806 3312 28858
rect 3336 28806 3346 28858
rect 3346 28806 3392 28858
rect 3416 28806 3462 28858
rect 3462 28806 3472 28858
rect 3496 28806 3526 28858
rect 3526 28806 3552 28858
rect 3256 28804 3312 28806
rect 3336 28804 3392 28806
rect 3416 28804 3472 28806
rect 3496 28804 3552 28806
rect 6256 28858 6312 28860
rect 6336 28858 6392 28860
rect 6416 28858 6472 28860
rect 6496 28858 6552 28860
rect 6256 28806 6282 28858
rect 6282 28806 6312 28858
rect 6336 28806 6346 28858
rect 6346 28806 6392 28858
rect 6416 28806 6462 28858
rect 6462 28806 6472 28858
rect 6496 28806 6526 28858
rect 6526 28806 6552 28858
rect 6256 28804 6312 28806
rect 6336 28804 6392 28806
rect 6416 28804 6472 28806
rect 6496 28804 6552 28806
rect 9256 28858 9312 28860
rect 9336 28858 9392 28860
rect 9416 28858 9472 28860
rect 9496 28858 9552 28860
rect 9256 28806 9282 28858
rect 9282 28806 9312 28858
rect 9336 28806 9346 28858
rect 9346 28806 9392 28858
rect 9416 28806 9462 28858
rect 9462 28806 9472 28858
rect 9496 28806 9526 28858
rect 9526 28806 9552 28858
rect 9256 28804 9312 28806
rect 9336 28804 9392 28806
rect 9416 28804 9472 28806
rect 9496 28804 9552 28806
rect 12256 28858 12312 28860
rect 12336 28858 12392 28860
rect 12416 28858 12472 28860
rect 12496 28858 12552 28860
rect 12256 28806 12282 28858
rect 12282 28806 12312 28858
rect 12336 28806 12346 28858
rect 12346 28806 12392 28858
rect 12416 28806 12462 28858
rect 12462 28806 12472 28858
rect 12496 28806 12526 28858
rect 12526 28806 12552 28858
rect 12256 28804 12312 28806
rect 12336 28804 12392 28806
rect 12416 28804 12472 28806
rect 12496 28804 12552 28806
rect 15256 28858 15312 28860
rect 15336 28858 15392 28860
rect 15416 28858 15472 28860
rect 15496 28858 15552 28860
rect 15256 28806 15282 28858
rect 15282 28806 15312 28858
rect 15336 28806 15346 28858
rect 15346 28806 15392 28858
rect 15416 28806 15462 28858
rect 15462 28806 15472 28858
rect 15496 28806 15526 28858
rect 15526 28806 15552 28858
rect 15256 28804 15312 28806
rect 15336 28804 15392 28806
rect 15416 28804 15472 28806
rect 15496 28804 15552 28806
rect 18256 28858 18312 28860
rect 18336 28858 18392 28860
rect 18416 28858 18472 28860
rect 18496 28858 18552 28860
rect 18256 28806 18282 28858
rect 18282 28806 18312 28858
rect 18336 28806 18346 28858
rect 18346 28806 18392 28858
rect 18416 28806 18462 28858
rect 18462 28806 18472 28858
rect 18496 28806 18526 28858
rect 18526 28806 18552 28858
rect 18256 28804 18312 28806
rect 18336 28804 18392 28806
rect 18416 28804 18472 28806
rect 18496 28804 18552 28806
rect 21256 28858 21312 28860
rect 21336 28858 21392 28860
rect 21416 28858 21472 28860
rect 21496 28858 21552 28860
rect 21256 28806 21282 28858
rect 21282 28806 21312 28858
rect 21336 28806 21346 28858
rect 21346 28806 21392 28858
rect 21416 28806 21462 28858
rect 21462 28806 21472 28858
rect 21496 28806 21526 28858
rect 21526 28806 21552 28858
rect 21256 28804 21312 28806
rect 21336 28804 21392 28806
rect 21416 28804 21472 28806
rect 21496 28804 21552 28806
rect 24256 28858 24312 28860
rect 24336 28858 24392 28860
rect 24416 28858 24472 28860
rect 24496 28858 24552 28860
rect 24256 28806 24282 28858
rect 24282 28806 24312 28858
rect 24336 28806 24346 28858
rect 24346 28806 24392 28858
rect 24416 28806 24462 28858
rect 24462 28806 24472 28858
rect 24496 28806 24526 28858
rect 24526 28806 24552 28858
rect 24256 28804 24312 28806
rect 24336 28804 24392 28806
rect 24416 28804 24472 28806
rect 24496 28804 24552 28806
rect 1756 28314 1812 28316
rect 1836 28314 1892 28316
rect 1916 28314 1972 28316
rect 1996 28314 2052 28316
rect 1756 28262 1782 28314
rect 1782 28262 1812 28314
rect 1836 28262 1846 28314
rect 1846 28262 1892 28314
rect 1916 28262 1962 28314
rect 1962 28262 1972 28314
rect 1996 28262 2026 28314
rect 2026 28262 2052 28314
rect 1756 28260 1812 28262
rect 1836 28260 1892 28262
rect 1916 28260 1972 28262
rect 1996 28260 2052 28262
rect 4756 28314 4812 28316
rect 4836 28314 4892 28316
rect 4916 28314 4972 28316
rect 4996 28314 5052 28316
rect 4756 28262 4782 28314
rect 4782 28262 4812 28314
rect 4836 28262 4846 28314
rect 4846 28262 4892 28314
rect 4916 28262 4962 28314
rect 4962 28262 4972 28314
rect 4996 28262 5026 28314
rect 5026 28262 5052 28314
rect 4756 28260 4812 28262
rect 4836 28260 4892 28262
rect 4916 28260 4972 28262
rect 4996 28260 5052 28262
rect 7756 28314 7812 28316
rect 7836 28314 7892 28316
rect 7916 28314 7972 28316
rect 7996 28314 8052 28316
rect 7756 28262 7782 28314
rect 7782 28262 7812 28314
rect 7836 28262 7846 28314
rect 7846 28262 7892 28314
rect 7916 28262 7962 28314
rect 7962 28262 7972 28314
rect 7996 28262 8026 28314
rect 8026 28262 8052 28314
rect 7756 28260 7812 28262
rect 7836 28260 7892 28262
rect 7916 28260 7972 28262
rect 7996 28260 8052 28262
rect 10756 28314 10812 28316
rect 10836 28314 10892 28316
rect 10916 28314 10972 28316
rect 10996 28314 11052 28316
rect 10756 28262 10782 28314
rect 10782 28262 10812 28314
rect 10836 28262 10846 28314
rect 10846 28262 10892 28314
rect 10916 28262 10962 28314
rect 10962 28262 10972 28314
rect 10996 28262 11026 28314
rect 11026 28262 11052 28314
rect 10756 28260 10812 28262
rect 10836 28260 10892 28262
rect 10916 28260 10972 28262
rect 10996 28260 11052 28262
rect 13756 28314 13812 28316
rect 13836 28314 13892 28316
rect 13916 28314 13972 28316
rect 13996 28314 14052 28316
rect 13756 28262 13782 28314
rect 13782 28262 13812 28314
rect 13836 28262 13846 28314
rect 13846 28262 13892 28314
rect 13916 28262 13962 28314
rect 13962 28262 13972 28314
rect 13996 28262 14026 28314
rect 14026 28262 14052 28314
rect 13756 28260 13812 28262
rect 13836 28260 13892 28262
rect 13916 28260 13972 28262
rect 13996 28260 14052 28262
rect 16756 28314 16812 28316
rect 16836 28314 16892 28316
rect 16916 28314 16972 28316
rect 16996 28314 17052 28316
rect 16756 28262 16782 28314
rect 16782 28262 16812 28314
rect 16836 28262 16846 28314
rect 16846 28262 16892 28314
rect 16916 28262 16962 28314
rect 16962 28262 16972 28314
rect 16996 28262 17026 28314
rect 17026 28262 17052 28314
rect 16756 28260 16812 28262
rect 16836 28260 16892 28262
rect 16916 28260 16972 28262
rect 16996 28260 17052 28262
rect 19756 28314 19812 28316
rect 19836 28314 19892 28316
rect 19916 28314 19972 28316
rect 19996 28314 20052 28316
rect 19756 28262 19782 28314
rect 19782 28262 19812 28314
rect 19836 28262 19846 28314
rect 19846 28262 19892 28314
rect 19916 28262 19962 28314
rect 19962 28262 19972 28314
rect 19996 28262 20026 28314
rect 20026 28262 20052 28314
rect 19756 28260 19812 28262
rect 19836 28260 19892 28262
rect 19916 28260 19972 28262
rect 19996 28260 20052 28262
rect 22756 28314 22812 28316
rect 22836 28314 22892 28316
rect 22916 28314 22972 28316
rect 22996 28314 23052 28316
rect 22756 28262 22782 28314
rect 22782 28262 22812 28314
rect 22836 28262 22846 28314
rect 22846 28262 22892 28314
rect 22916 28262 22962 28314
rect 22962 28262 22972 28314
rect 22996 28262 23026 28314
rect 23026 28262 23052 28314
rect 22756 28260 22812 28262
rect 22836 28260 22892 28262
rect 22916 28260 22972 28262
rect 22996 28260 23052 28262
rect 3256 27770 3312 27772
rect 3336 27770 3392 27772
rect 3416 27770 3472 27772
rect 3496 27770 3552 27772
rect 3256 27718 3282 27770
rect 3282 27718 3312 27770
rect 3336 27718 3346 27770
rect 3346 27718 3392 27770
rect 3416 27718 3462 27770
rect 3462 27718 3472 27770
rect 3496 27718 3526 27770
rect 3526 27718 3552 27770
rect 3256 27716 3312 27718
rect 3336 27716 3392 27718
rect 3416 27716 3472 27718
rect 3496 27716 3552 27718
rect 6256 27770 6312 27772
rect 6336 27770 6392 27772
rect 6416 27770 6472 27772
rect 6496 27770 6552 27772
rect 6256 27718 6282 27770
rect 6282 27718 6312 27770
rect 6336 27718 6346 27770
rect 6346 27718 6392 27770
rect 6416 27718 6462 27770
rect 6462 27718 6472 27770
rect 6496 27718 6526 27770
rect 6526 27718 6552 27770
rect 6256 27716 6312 27718
rect 6336 27716 6392 27718
rect 6416 27716 6472 27718
rect 6496 27716 6552 27718
rect 9256 27770 9312 27772
rect 9336 27770 9392 27772
rect 9416 27770 9472 27772
rect 9496 27770 9552 27772
rect 9256 27718 9282 27770
rect 9282 27718 9312 27770
rect 9336 27718 9346 27770
rect 9346 27718 9392 27770
rect 9416 27718 9462 27770
rect 9462 27718 9472 27770
rect 9496 27718 9526 27770
rect 9526 27718 9552 27770
rect 9256 27716 9312 27718
rect 9336 27716 9392 27718
rect 9416 27716 9472 27718
rect 9496 27716 9552 27718
rect 12256 27770 12312 27772
rect 12336 27770 12392 27772
rect 12416 27770 12472 27772
rect 12496 27770 12552 27772
rect 12256 27718 12282 27770
rect 12282 27718 12312 27770
rect 12336 27718 12346 27770
rect 12346 27718 12392 27770
rect 12416 27718 12462 27770
rect 12462 27718 12472 27770
rect 12496 27718 12526 27770
rect 12526 27718 12552 27770
rect 12256 27716 12312 27718
rect 12336 27716 12392 27718
rect 12416 27716 12472 27718
rect 12496 27716 12552 27718
rect 15256 27770 15312 27772
rect 15336 27770 15392 27772
rect 15416 27770 15472 27772
rect 15496 27770 15552 27772
rect 15256 27718 15282 27770
rect 15282 27718 15312 27770
rect 15336 27718 15346 27770
rect 15346 27718 15392 27770
rect 15416 27718 15462 27770
rect 15462 27718 15472 27770
rect 15496 27718 15526 27770
rect 15526 27718 15552 27770
rect 15256 27716 15312 27718
rect 15336 27716 15392 27718
rect 15416 27716 15472 27718
rect 15496 27716 15552 27718
rect 18256 27770 18312 27772
rect 18336 27770 18392 27772
rect 18416 27770 18472 27772
rect 18496 27770 18552 27772
rect 18256 27718 18282 27770
rect 18282 27718 18312 27770
rect 18336 27718 18346 27770
rect 18346 27718 18392 27770
rect 18416 27718 18462 27770
rect 18462 27718 18472 27770
rect 18496 27718 18526 27770
rect 18526 27718 18552 27770
rect 18256 27716 18312 27718
rect 18336 27716 18392 27718
rect 18416 27716 18472 27718
rect 18496 27716 18552 27718
rect 21256 27770 21312 27772
rect 21336 27770 21392 27772
rect 21416 27770 21472 27772
rect 21496 27770 21552 27772
rect 21256 27718 21282 27770
rect 21282 27718 21312 27770
rect 21336 27718 21346 27770
rect 21346 27718 21392 27770
rect 21416 27718 21462 27770
rect 21462 27718 21472 27770
rect 21496 27718 21526 27770
rect 21526 27718 21552 27770
rect 21256 27716 21312 27718
rect 21336 27716 21392 27718
rect 21416 27716 21472 27718
rect 21496 27716 21552 27718
rect 24256 27770 24312 27772
rect 24336 27770 24392 27772
rect 24416 27770 24472 27772
rect 24496 27770 24552 27772
rect 24256 27718 24282 27770
rect 24282 27718 24312 27770
rect 24336 27718 24346 27770
rect 24346 27718 24392 27770
rect 24416 27718 24462 27770
rect 24462 27718 24472 27770
rect 24496 27718 24526 27770
rect 24526 27718 24552 27770
rect 24256 27716 24312 27718
rect 24336 27716 24392 27718
rect 24416 27716 24472 27718
rect 24496 27716 24552 27718
rect 25756 29402 25812 29404
rect 25836 29402 25892 29404
rect 25916 29402 25972 29404
rect 25996 29402 26052 29404
rect 25756 29350 25782 29402
rect 25782 29350 25812 29402
rect 25836 29350 25846 29402
rect 25846 29350 25892 29402
rect 25916 29350 25962 29402
rect 25962 29350 25972 29402
rect 25996 29350 26026 29402
rect 26026 29350 26052 29402
rect 25756 29348 25812 29350
rect 25836 29348 25892 29350
rect 25916 29348 25972 29350
rect 25996 29348 26052 29350
rect 27256 28858 27312 28860
rect 27336 28858 27392 28860
rect 27416 28858 27472 28860
rect 27496 28858 27552 28860
rect 27256 28806 27282 28858
rect 27282 28806 27312 28858
rect 27336 28806 27346 28858
rect 27346 28806 27392 28858
rect 27416 28806 27462 28858
rect 27462 28806 27472 28858
rect 27496 28806 27526 28858
rect 27526 28806 27552 28858
rect 27256 28804 27312 28806
rect 27336 28804 27392 28806
rect 27416 28804 27472 28806
rect 27496 28804 27552 28806
rect 25756 28314 25812 28316
rect 25836 28314 25892 28316
rect 25916 28314 25972 28316
rect 25996 28314 26052 28316
rect 25756 28262 25782 28314
rect 25782 28262 25812 28314
rect 25836 28262 25846 28314
rect 25846 28262 25892 28314
rect 25916 28262 25962 28314
rect 25962 28262 25972 28314
rect 25996 28262 26026 28314
rect 26026 28262 26052 28314
rect 25756 28260 25812 28262
rect 25836 28260 25892 28262
rect 25916 28260 25972 28262
rect 25996 28260 26052 28262
rect 27256 27770 27312 27772
rect 27336 27770 27392 27772
rect 27416 27770 27472 27772
rect 27496 27770 27552 27772
rect 27256 27718 27282 27770
rect 27282 27718 27312 27770
rect 27336 27718 27346 27770
rect 27346 27718 27392 27770
rect 27416 27718 27462 27770
rect 27462 27718 27472 27770
rect 27496 27718 27526 27770
rect 27526 27718 27552 27770
rect 27256 27716 27312 27718
rect 27336 27716 27392 27718
rect 27416 27716 27472 27718
rect 27496 27716 27552 27718
rect 1756 27226 1812 27228
rect 1836 27226 1892 27228
rect 1916 27226 1972 27228
rect 1996 27226 2052 27228
rect 1756 27174 1782 27226
rect 1782 27174 1812 27226
rect 1836 27174 1846 27226
rect 1846 27174 1892 27226
rect 1916 27174 1962 27226
rect 1962 27174 1972 27226
rect 1996 27174 2026 27226
rect 2026 27174 2052 27226
rect 1756 27172 1812 27174
rect 1836 27172 1892 27174
rect 1916 27172 1972 27174
rect 1996 27172 2052 27174
rect 4756 27226 4812 27228
rect 4836 27226 4892 27228
rect 4916 27226 4972 27228
rect 4996 27226 5052 27228
rect 4756 27174 4782 27226
rect 4782 27174 4812 27226
rect 4836 27174 4846 27226
rect 4846 27174 4892 27226
rect 4916 27174 4962 27226
rect 4962 27174 4972 27226
rect 4996 27174 5026 27226
rect 5026 27174 5052 27226
rect 4756 27172 4812 27174
rect 4836 27172 4892 27174
rect 4916 27172 4972 27174
rect 4996 27172 5052 27174
rect 7756 27226 7812 27228
rect 7836 27226 7892 27228
rect 7916 27226 7972 27228
rect 7996 27226 8052 27228
rect 7756 27174 7782 27226
rect 7782 27174 7812 27226
rect 7836 27174 7846 27226
rect 7846 27174 7892 27226
rect 7916 27174 7962 27226
rect 7962 27174 7972 27226
rect 7996 27174 8026 27226
rect 8026 27174 8052 27226
rect 7756 27172 7812 27174
rect 7836 27172 7892 27174
rect 7916 27172 7972 27174
rect 7996 27172 8052 27174
rect 10756 27226 10812 27228
rect 10836 27226 10892 27228
rect 10916 27226 10972 27228
rect 10996 27226 11052 27228
rect 10756 27174 10782 27226
rect 10782 27174 10812 27226
rect 10836 27174 10846 27226
rect 10846 27174 10892 27226
rect 10916 27174 10962 27226
rect 10962 27174 10972 27226
rect 10996 27174 11026 27226
rect 11026 27174 11052 27226
rect 10756 27172 10812 27174
rect 10836 27172 10892 27174
rect 10916 27172 10972 27174
rect 10996 27172 11052 27174
rect 13756 27226 13812 27228
rect 13836 27226 13892 27228
rect 13916 27226 13972 27228
rect 13996 27226 14052 27228
rect 13756 27174 13782 27226
rect 13782 27174 13812 27226
rect 13836 27174 13846 27226
rect 13846 27174 13892 27226
rect 13916 27174 13962 27226
rect 13962 27174 13972 27226
rect 13996 27174 14026 27226
rect 14026 27174 14052 27226
rect 13756 27172 13812 27174
rect 13836 27172 13892 27174
rect 13916 27172 13972 27174
rect 13996 27172 14052 27174
rect 16756 27226 16812 27228
rect 16836 27226 16892 27228
rect 16916 27226 16972 27228
rect 16996 27226 17052 27228
rect 16756 27174 16782 27226
rect 16782 27174 16812 27226
rect 16836 27174 16846 27226
rect 16846 27174 16892 27226
rect 16916 27174 16962 27226
rect 16962 27174 16972 27226
rect 16996 27174 17026 27226
rect 17026 27174 17052 27226
rect 16756 27172 16812 27174
rect 16836 27172 16892 27174
rect 16916 27172 16972 27174
rect 16996 27172 17052 27174
rect 19756 27226 19812 27228
rect 19836 27226 19892 27228
rect 19916 27226 19972 27228
rect 19996 27226 20052 27228
rect 19756 27174 19782 27226
rect 19782 27174 19812 27226
rect 19836 27174 19846 27226
rect 19846 27174 19892 27226
rect 19916 27174 19962 27226
rect 19962 27174 19972 27226
rect 19996 27174 20026 27226
rect 20026 27174 20052 27226
rect 19756 27172 19812 27174
rect 19836 27172 19892 27174
rect 19916 27172 19972 27174
rect 19996 27172 20052 27174
rect 22756 27226 22812 27228
rect 22836 27226 22892 27228
rect 22916 27226 22972 27228
rect 22996 27226 23052 27228
rect 22756 27174 22782 27226
rect 22782 27174 22812 27226
rect 22836 27174 22846 27226
rect 22846 27174 22892 27226
rect 22916 27174 22962 27226
rect 22962 27174 22972 27226
rect 22996 27174 23026 27226
rect 23026 27174 23052 27226
rect 22756 27172 22812 27174
rect 22836 27172 22892 27174
rect 22916 27172 22972 27174
rect 22996 27172 23052 27174
rect 3256 26682 3312 26684
rect 3336 26682 3392 26684
rect 3416 26682 3472 26684
rect 3496 26682 3552 26684
rect 3256 26630 3282 26682
rect 3282 26630 3312 26682
rect 3336 26630 3346 26682
rect 3346 26630 3392 26682
rect 3416 26630 3462 26682
rect 3462 26630 3472 26682
rect 3496 26630 3526 26682
rect 3526 26630 3552 26682
rect 3256 26628 3312 26630
rect 3336 26628 3392 26630
rect 3416 26628 3472 26630
rect 3496 26628 3552 26630
rect 6256 26682 6312 26684
rect 6336 26682 6392 26684
rect 6416 26682 6472 26684
rect 6496 26682 6552 26684
rect 6256 26630 6282 26682
rect 6282 26630 6312 26682
rect 6336 26630 6346 26682
rect 6346 26630 6392 26682
rect 6416 26630 6462 26682
rect 6462 26630 6472 26682
rect 6496 26630 6526 26682
rect 6526 26630 6552 26682
rect 6256 26628 6312 26630
rect 6336 26628 6392 26630
rect 6416 26628 6472 26630
rect 6496 26628 6552 26630
rect 9256 26682 9312 26684
rect 9336 26682 9392 26684
rect 9416 26682 9472 26684
rect 9496 26682 9552 26684
rect 9256 26630 9282 26682
rect 9282 26630 9312 26682
rect 9336 26630 9346 26682
rect 9346 26630 9392 26682
rect 9416 26630 9462 26682
rect 9462 26630 9472 26682
rect 9496 26630 9526 26682
rect 9526 26630 9552 26682
rect 9256 26628 9312 26630
rect 9336 26628 9392 26630
rect 9416 26628 9472 26630
rect 9496 26628 9552 26630
rect 12256 26682 12312 26684
rect 12336 26682 12392 26684
rect 12416 26682 12472 26684
rect 12496 26682 12552 26684
rect 12256 26630 12282 26682
rect 12282 26630 12312 26682
rect 12336 26630 12346 26682
rect 12346 26630 12392 26682
rect 12416 26630 12462 26682
rect 12462 26630 12472 26682
rect 12496 26630 12526 26682
rect 12526 26630 12552 26682
rect 12256 26628 12312 26630
rect 12336 26628 12392 26630
rect 12416 26628 12472 26630
rect 12496 26628 12552 26630
rect 15256 26682 15312 26684
rect 15336 26682 15392 26684
rect 15416 26682 15472 26684
rect 15496 26682 15552 26684
rect 15256 26630 15282 26682
rect 15282 26630 15312 26682
rect 15336 26630 15346 26682
rect 15346 26630 15392 26682
rect 15416 26630 15462 26682
rect 15462 26630 15472 26682
rect 15496 26630 15526 26682
rect 15526 26630 15552 26682
rect 15256 26628 15312 26630
rect 15336 26628 15392 26630
rect 15416 26628 15472 26630
rect 15496 26628 15552 26630
rect 18256 26682 18312 26684
rect 18336 26682 18392 26684
rect 18416 26682 18472 26684
rect 18496 26682 18552 26684
rect 18256 26630 18282 26682
rect 18282 26630 18312 26682
rect 18336 26630 18346 26682
rect 18346 26630 18392 26682
rect 18416 26630 18462 26682
rect 18462 26630 18472 26682
rect 18496 26630 18526 26682
rect 18526 26630 18552 26682
rect 18256 26628 18312 26630
rect 18336 26628 18392 26630
rect 18416 26628 18472 26630
rect 18496 26628 18552 26630
rect 21256 26682 21312 26684
rect 21336 26682 21392 26684
rect 21416 26682 21472 26684
rect 21496 26682 21552 26684
rect 21256 26630 21282 26682
rect 21282 26630 21312 26682
rect 21336 26630 21346 26682
rect 21346 26630 21392 26682
rect 21416 26630 21462 26682
rect 21462 26630 21472 26682
rect 21496 26630 21526 26682
rect 21526 26630 21552 26682
rect 21256 26628 21312 26630
rect 21336 26628 21392 26630
rect 21416 26628 21472 26630
rect 21496 26628 21552 26630
rect 1756 26138 1812 26140
rect 1836 26138 1892 26140
rect 1916 26138 1972 26140
rect 1996 26138 2052 26140
rect 1756 26086 1782 26138
rect 1782 26086 1812 26138
rect 1836 26086 1846 26138
rect 1846 26086 1892 26138
rect 1916 26086 1962 26138
rect 1962 26086 1972 26138
rect 1996 26086 2026 26138
rect 2026 26086 2052 26138
rect 1756 26084 1812 26086
rect 1836 26084 1892 26086
rect 1916 26084 1972 26086
rect 1996 26084 2052 26086
rect 4756 26138 4812 26140
rect 4836 26138 4892 26140
rect 4916 26138 4972 26140
rect 4996 26138 5052 26140
rect 4756 26086 4782 26138
rect 4782 26086 4812 26138
rect 4836 26086 4846 26138
rect 4846 26086 4892 26138
rect 4916 26086 4962 26138
rect 4962 26086 4972 26138
rect 4996 26086 5026 26138
rect 5026 26086 5052 26138
rect 4756 26084 4812 26086
rect 4836 26084 4892 26086
rect 4916 26084 4972 26086
rect 4996 26084 5052 26086
rect 7756 26138 7812 26140
rect 7836 26138 7892 26140
rect 7916 26138 7972 26140
rect 7996 26138 8052 26140
rect 7756 26086 7782 26138
rect 7782 26086 7812 26138
rect 7836 26086 7846 26138
rect 7846 26086 7892 26138
rect 7916 26086 7962 26138
rect 7962 26086 7972 26138
rect 7996 26086 8026 26138
rect 8026 26086 8052 26138
rect 7756 26084 7812 26086
rect 7836 26084 7892 26086
rect 7916 26084 7972 26086
rect 7996 26084 8052 26086
rect 10756 26138 10812 26140
rect 10836 26138 10892 26140
rect 10916 26138 10972 26140
rect 10996 26138 11052 26140
rect 10756 26086 10782 26138
rect 10782 26086 10812 26138
rect 10836 26086 10846 26138
rect 10846 26086 10892 26138
rect 10916 26086 10962 26138
rect 10962 26086 10972 26138
rect 10996 26086 11026 26138
rect 11026 26086 11052 26138
rect 10756 26084 10812 26086
rect 10836 26084 10892 26086
rect 10916 26084 10972 26086
rect 10996 26084 11052 26086
rect 13756 26138 13812 26140
rect 13836 26138 13892 26140
rect 13916 26138 13972 26140
rect 13996 26138 14052 26140
rect 13756 26086 13782 26138
rect 13782 26086 13812 26138
rect 13836 26086 13846 26138
rect 13846 26086 13892 26138
rect 13916 26086 13962 26138
rect 13962 26086 13972 26138
rect 13996 26086 14026 26138
rect 14026 26086 14052 26138
rect 13756 26084 13812 26086
rect 13836 26084 13892 26086
rect 13916 26084 13972 26086
rect 13996 26084 14052 26086
rect 16756 26138 16812 26140
rect 16836 26138 16892 26140
rect 16916 26138 16972 26140
rect 16996 26138 17052 26140
rect 16756 26086 16782 26138
rect 16782 26086 16812 26138
rect 16836 26086 16846 26138
rect 16846 26086 16892 26138
rect 16916 26086 16962 26138
rect 16962 26086 16972 26138
rect 16996 26086 17026 26138
rect 17026 26086 17052 26138
rect 16756 26084 16812 26086
rect 16836 26084 16892 26086
rect 16916 26084 16972 26086
rect 16996 26084 17052 26086
rect 19756 26138 19812 26140
rect 19836 26138 19892 26140
rect 19916 26138 19972 26140
rect 19996 26138 20052 26140
rect 19756 26086 19782 26138
rect 19782 26086 19812 26138
rect 19836 26086 19846 26138
rect 19846 26086 19892 26138
rect 19916 26086 19962 26138
rect 19962 26086 19972 26138
rect 19996 26086 20026 26138
rect 20026 26086 20052 26138
rect 19756 26084 19812 26086
rect 19836 26084 19892 26086
rect 19916 26084 19972 26086
rect 19996 26084 20052 26086
rect 22756 26138 22812 26140
rect 22836 26138 22892 26140
rect 22916 26138 22972 26140
rect 22996 26138 23052 26140
rect 22756 26086 22782 26138
rect 22782 26086 22812 26138
rect 22836 26086 22846 26138
rect 22846 26086 22892 26138
rect 22916 26086 22962 26138
rect 22962 26086 22972 26138
rect 22996 26086 23026 26138
rect 23026 26086 23052 26138
rect 22756 26084 22812 26086
rect 22836 26084 22892 26086
rect 22916 26084 22972 26086
rect 22996 26084 23052 26086
rect 3256 25594 3312 25596
rect 3336 25594 3392 25596
rect 3416 25594 3472 25596
rect 3496 25594 3552 25596
rect 3256 25542 3282 25594
rect 3282 25542 3312 25594
rect 3336 25542 3346 25594
rect 3346 25542 3392 25594
rect 3416 25542 3462 25594
rect 3462 25542 3472 25594
rect 3496 25542 3526 25594
rect 3526 25542 3552 25594
rect 3256 25540 3312 25542
rect 3336 25540 3392 25542
rect 3416 25540 3472 25542
rect 3496 25540 3552 25542
rect 6256 25594 6312 25596
rect 6336 25594 6392 25596
rect 6416 25594 6472 25596
rect 6496 25594 6552 25596
rect 6256 25542 6282 25594
rect 6282 25542 6312 25594
rect 6336 25542 6346 25594
rect 6346 25542 6392 25594
rect 6416 25542 6462 25594
rect 6462 25542 6472 25594
rect 6496 25542 6526 25594
rect 6526 25542 6552 25594
rect 6256 25540 6312 25542
rect 6336 25540 6392 25542
rect 6416 25540 6472 25542
rect 6496 25540 6552 25542
rect 9256 25594 9312 25596
rect 9336 25594 9392 25596
rect 9416 25594 9472 25596
rect 9496 25594 9552 25596
rect 9256 25542 9282 25594
rect 9282 25542 9312 25594
rect 9336 25542 9346 25594
rect 9346 25542 9392 25594
rect 9416 25542 9462 25594
rect 9462 25542 9472 25594
rect 9496 25542 9526 25594
rect 9526 25542 9552 25594
rect 9256 25540 9312 25542
rect 9336 25540 9392 25542
rect 9416 25540 9472 25542
rect 9496 25540 9552 25542
rect 12256 25594 12312 25596
rect 12336 25594 12392 25596
rect 12416 25594 12472 25596
rect 12496 25594 12552 25596
rect 12256 25542 12282 25594
rect 12282 25542 12312 25594
rect 12336 25542 12346 25594
rect 12346 25542 12392 25594
rect 12416 25542 12462 25594
rect 12462 25542 12472 25594
rect 12496 25542 12526 25594
rect 12526 25542 12552 25594
rect 12256 25540 12312 25542
rect 12336 25540 12392 25542
rect 12416 25540 12472 25542
rect 12496 25540 12552 25542
rect 15256 25594 15312 25596
rect 15336 25594 15392 25596
rect 15416 25594 15472 25596
rect 15496 25594 15552 25596
rect 15256 25542 15282 25594
rect 15282 25542 15312 25594
rect 15336 25542 15346 25594
rect 15346 25542 15392 25594
rect 15416 25542 15462 25594
rect 15462 25542 15472 25594
rect 15496 25542 15526 25594
rect 15526 25542 15552 25594
rect 15256 25540 15312 25542
rect 15336 25540 15392 25542
rect 15416 25540 15472 25542
rect 15496 25540 15552 25542
rect 18256 25594 18312 25596
rect 18336 25594 18392 25596
rect 18416 25594 18472 25596
rect 18496 25594 18552 25596
rect 18256 25542 18282 25594
rect 18282 25542 18312 25594
rect 18336 25542 18346 25594
rect 18346 25542 18392 25594
rect 18416 25542 18462 25594
rect 18462 25542 18472 25594
rect 18496 25542 18526 25594
rect 18526 25542 18552 25594
rect 18256 25540 18312 25542
rect 18336 25540 18392 25542
rect 18416 25540 18472 25542
rect 18496 25540 18552 25542
rect 21256 25594 21312 25596
rect 21336 25594 21392 25596
rect 21416 25594 21472 25596
rect 21496 25594 21552 25596
rect 21256 25542 21282 25594
rect 21282 25542 21312 25594
rect 21336 25542 21346 25594
rect 21346 25542 21392 25594
rect 21416 25542 21462 25594
rect 21462 25542 21472 25594
rect 21496 25542 21526 25594
rect 21526 25542 21552 25594
rect 21256 25540 21312 25542
rect 21336 25540 21392 25542
rect 21416 25540 21472 25542
rect 21496 25540 21552 25542
rect 1756 25050 1812 25052
rect 1836 25050 1892 25052
rect 1916 25050 1972 25052
rect 1996 25050 2052 25052
rect 1756 24998 1782 25050
rect 1782 24998 1812 25050
rect 1836 24998 1846 25050
rect 1846 24998 1892 25050
rect 1916 24998 1962 25050
rect 1962 24998 1972 25050
rect 1996 24998 2026 25050
rect 2026 24998 2052 25050
rect 1756 24996 1812 24998
rect 1836 24996 1892 24998
rect 1916 24996 1972 24998
rect 1996 24996 2052 24998
rect 4756 25050 4812 25052
rect 4836 25050 4892 25052
rect 4916 25050 4972 25052
rect 4996 25050 5052 25052
rect 4756 24998 4782 25050
rect 4782 24998 4812 25050
rect 4836 24998 4846 25050
rect 4846 24998 4892 25050
rect 4916 24998 4962 25050
rect 4962 24998 4972 25050
rect 4996 24998 5026 25050
rect 5026 24998 5052 25050
rect 4756 24996 4812 24998
rect 4836 24996 4892 24998
rect 4916 24996 4972 24998
rect 4996 24996 5052 24998
rect 7756 25050 7812 25052
rect 7836 25050 7892 25052
rect 7916 25050 7972 25052
rect 7996 25050 8052 25052
rect 7756 24998 7782 25050
rect 7782 24998 7812 25050
rect 7836 24998 7846 25050
rect 7846 24998 7892 25050
rect 7916 24998 7962 25050
rect 7962 24998 7972 25050
rect 7996 24998 8026 25050
rect 8026 24998 8052 25050
rect 7756 24996 7812 24998
rect 7836 24996 7892 24998
rect 7916 24996 7972 24998
rect 7996 24996 8052 24998
rect 10756 25050 10812 25052
rect 10836 25050 10892 25052
rect 10916 25050 10972 25052
rect 10996 25050 11052 25052
rect 10756 24998 10782 25050
rect 10782 24998 10812 25050
rect 10836 24998 10846 25050
rect 10846 24998 10892 25050
rect 10916 24998 10962 25050
rect 10962 24998 10972 25050
rect 10996 24998 11026 25050
rect 11026 24998 11052 25050
rect 10756 24996 10812 24998
rect 10836 24996 10892 24998
rect 10916 24996 10972 24998
rect 10996 24996 11052 24998
rect 13756 25050 13812 25052
rect 13836 25050 13892 25052
rect 13916 25050 13972 25052
rect 13996 25050 14052 25052
rect 13756 24998 13782 25050
rect 13782 24998 13812 25050
rect 13836 24998 13846 25050
rect 13846 24998 13892 25050
rect 13916 24998 13962 25050
rect 13962 24998 13972 25050
rect 13996 24998 14026 25050
rect 14026 24998 14052 25050
rect 13756 24996 13812 24998
rect 13836 24996 13892 24998
rect 13916 24996 13972 24998
rect 13996 24996 14052 24998
rect 16756 25050 16812 25052
rect 16836 25050 16892 25052
rect 16916 25050 16972 25052
rect 16996 25050 17052 25052
rect 16756 24998 16782 25050
rect 16782 24998 16812 25050
rect 16836 24998 16846 25050
rect 16846 24998 16892 25050
rect 16916 24998 16962 25050
rect 16962 24998 16972 25050
rect 16996 24998 17026 25050
rect 17026 24998 17052 25050
rect 16756 24996 16812 24998
rect 16836 24996 16892 24998
rect 16916 24996 16972 24998
rect 16996 24996 17052 24998
rect 19756 25050 19812 25052
rect 19836 25050 19892 25052
rect 19916 25050 19972 25052
rect 19996 25050 20052 25052
rect 19756 24998 19782 25050
rect 19782 24998 19812 25050
rect 19836 24998 19846 25050
rect 19846 24998 19892 25050
rect 19916 24998 19962 25050
rect 19962 24998 19972 25050
rect 19996 24998 20026 25050
rect 20026 24998 20052 25050
rect 19756 24996 19812 24998
rect 19836 24996 19892 24998
rect 19916 24996 19972 24998
rect 19996 24996 20052 24998
rect 22756 25050 22812 25052
rect 22836 25050 22892 25052
rect 22916 25050 22972 25052
rect 22996 25050 23052 25052
rect 22756 24998 22782 25050
rect 22782 24998 22812 25050
rect 22836 24998 22846 25050
rect 22846 24998 22892 25050
rect 22916 24998 22962 25050
rect 22962 24998 22972 25050
rect 22996 24998 23026 25050
rect 23026 24998 23052 25050
rect 22756 24996 22812 24998
rect 22836 24996 22892 24998
rect 22916 24996 22972 24998
rect 22996 24996 23052 24998
rect 3256 24506 3312 24508
rect 3336 24506 3392 24508
rect 3416 24506 3472 24508
rect 3496 24506 3552 24508
rect 3256 24454 3282 24506
rect 3282 24454 3312 24506
rect 3336 24454 3346 24506
rect 3346 24454 3392 24506
rect 3416 24454 3462 24506
rect 3462 24454 3472 24506
rect 3496 24454 3526 24506
rect 3526 24454 3552 24506
rect 3256 24452 3312 24454
rect 3336 24452 3392 24454
rect 3416 24452 3472 24454
rect 3496 24452 3552 24454
rect 6256 24506 6312 24508
rect 6336 24506 6392 24508
rect 6416 24506 6472 24508
rect 6496 24506 6552 24508
rect 6256 24454 6282 24506
rect 6282 24454 6312 24506
rect 6336 24454 6346 24506
rect 6346 24454 6392 24506
rect 6416 24454 6462 24506
rect 6462 24454 6472 24506
rect 6496 24454 6526 24506
rect 6526 24454 6552 24506
rect 6256 24452 6312 24454
rect 6336 24452 6392 24454
rect 6416 24452 6472 24454
rect 6496 24452 6552 24454
rect 9256 24506 9312 24508
rect 9336 24506 9392 24508
rect 9416 24506 9472 24508
rect 9496 24506 9552 24508
rect 9256 24454 9282 24506
rect 9282 24454 9312 24506
rect 9336 24454 9346 24506
rect 9346 24454 9392 24506
rect 9416 24454 9462 24506
rect 9462 24454 9472 24506
rect 9496 24454 9526 24506
rect 9526 24454 9552 24506
rect 9256 24452 9312 24454
rect 9336 24452 9392 24454
rect 9416 24452 9472 24454
rect 9496 24452 9552 24454
rect 12256 24506 12312 24508
rect 12336 24506 12392 24508
rect 12416 24506 12472 24508
rect 12496 24506 12552 24508
rect 12256 24454 12282 24506
rect 12282 24454 12312 24506
rect 12336 24454 12346 24506
rect 12346 24454 12392 24506
rect 12416 24454 12462 24506
rect 12462 24454 12472 24506
rect 12496 24454 12526 24506
rect 12526 24454 12552 24506
rect 12256 24452 12312 24454
rect 12336 24452 12392 24454
rect 12416 24452 12472 24454
rect 12496 24452 12552 24454
rect 15256 24506 15312 24508
rect 15336 24506 15392 24508
rect 15416 24506 15472 24508
rect 15496 24506 15552 24508
rect 15256 24454 15282 24506
rect 15282 24454 15312 24506
rect 15336 24454 15346 24506
rect 15346 24454 15392 24506
rect 15416 24454 15462 24506
rect 15462 24454 15472 24506
rect 15496 24454 15526 24506
rect 15526 24454 15552 24506
rect 15256 24452 15312 24454
rect 15336 24452 15392 24454
rect 15416 24452 15472 24454
rect 15496 24452 15552 24454
rect 18256 24506 18312 24508
rect 18336 24506 18392 24508
rect 18416 24506 18472 24508
rect 18496 24506 18552 24508
rect 18256 24454 18282 24506
rect 18282 24454 18312 24506
rect 18336 24454 18346 24506
rect 18346 24454 18392 24506
rect 18416 24454 18462 24506
rect 18462 24454 18472 24506
rect 18496 24454 18526 24506
rect 18526 24454 18552 24506
rect 18256 24452 18312 24454
rect 18336 24452 18392 24454
rect 18416 24452 18472 24454
rect 18496 24452 18552 24454
rect 21256 24506 21312 24508
rect 21336 24506 21392 24508
rect 21416 24506 21472 24508
rect 21496 24506 21552 24508
rect 21256 24454 21282 24506
rect 21282 24454 21312 24506
rect 21336 24454 21346 24506
rect 21346 24454 21392 24506
rect 21416 24454 21462 24506
rect 21462 24454 21472 24506
rect 21496 24454 21526 24506
rect 21526 24454 21552 24506
rect 21256 24452 21312 24454
rect 21336 24452 21392 24454
rect 21416 24452 21472 24454
rect 21496 24452 21552 24454
rect 1756 23962 1812 23964
rect 1836 23962 1892 23964
rect 1916 23962 1972 23964
rect 1996 23962 2052 23964
rect 1756 23910 1782 23962
rect 1782 23910 1812 23962
rect 1836 23910 1846 23962
rect 1846 23910 1892 23962
rect 1916 23910 1962 23962
rect 1962 23910 1972 23962
rect 1996 23910 2026 23962
rect 2026 23910 2052 23962
rect 1756 23908 1812 23910
rect 1836 23908 1892 23910
rect 1916 23908 1972 23910
rect 1996 23908 2052 23910
rect 4756 23962 4812 23964
rect 4836 23962 4892 23964
rect 4916 23962 4972 23964
rect 4996 23962 5052 23964
rect 4756 23910 4782 23962
rect 4782 23910 4812 23962
rect 4836 23910 4846 23962
rect 4846 23910 4892 23962
rect 4916 23910 4962 23962
rect 4962 23910 4972 23962
rect 4996 23910 5026 23962
rect 5026 23910 5052 23962
rect 4756 23908 4812 23910
rect 4836 23908 4892 23910
rect 4916 23908 4972 23910
rect 4996 23908 5052 23910
rect 7756 23962 7812 23964
rect 7836 23962 7892 23964
rect 7916 23962 7972 23964
rect 7996 23962 8052 23964
rect 7756 23910 7782 23962
rect 7782 23910 7812 23962
rect 7836 23910 7846 23962
rect 7846 23910 7892 23962
rect 7916 23910 7962 23962
rect 7962 23910 7972 23962
rect 7996 23910 8026 23962
rect 8026 23910 8052 23962
rect 7756 23908 7812 23910
rect 7836 23908 7892 23910
rect 7916 23908 7972 23910
rect 7996 23908 8052 23910
rect 10756 23962 10812 23964
rect 10836 23962 10892 23964
rect 10916 23962 10972 23964
rect 10996 23962 11052 23964
rect 10756 23910 10782 23962
rect 10782 23910 10812 23962
rect 10836 23910 10846 23962
rect 10846 23910 10892 23962
rect 10916 23910 10962 23962
rect 10962 23910 10972 23962
rect 10996 23910 11026 23962
rect 11026 23910 11052 23962
rect 10756 23908 10812 23910
rect 10836 23908 10892 23910
rect 10916 23908 10972 23910
rect 10996 23908 11052 23910
rect 13756 23962 13812 23964
rect 13836 23962 13892 23964
rect 13916 23962 13972 23964
rect 13996 23962 14052 23964
rect 13756 23910 13782 23962
rect 13782 23910 13812 23962
rect 13836 23910 13846 23962
rect 13846 23910 13892 23962
rect 13916 23910 13962 23962
rect 13962 23910 13972 23962
rect 13996 23910 14026 23962
rect 14026 23910 14052 23962
rect 13756 23908 13812 23910
rect 13836 23908 13892 23910
rect 13916 23908 13972 23910
rect 13996 23908 14052 23910
rect 16756 23962 16812 23964
rect 16836 23962 16892 23964
rect 16916 23962 16972 23964
rect 16996 23962 17052 23964
rect 16756 23910 16782 23962
rect 16782 23910 16812 23962
rect 16836 23910 16846 23962
rect 16846 23910 16892 23962
rect 16916 23910 16962 23962
rect 16962 23910 16972 23962
rect 16996 23910 17026 23962
rect 17026 23910 17052 23962
rect 16756 23908 16812 23910
rect 16836 23908 16892 23910
rect 16916 23908 16972 23910
rect 16996 23908 17052 23910
rect 19756 23962 19812 23964
rect 19836 23962 19892 23964
rect 19916 23962 19972 23964
rect 19996 23962 20052 23964
rect 19756 23910 19782 23962
rect 19782 23910 19812 23962
rect 19836 23910 19846 23962
rect 19846 23910 19892 23962
rect 19916 23910 19962 23962
rect 19962 23910 19972 23962
rect 19996 23910 20026 23962
rect 20026 23910 20052 23962
rect 19756 23908 19812 23910
rect 19836 23908 19892 23910
rect 19916 23908 19972 23910
rect 19996 23908 20052 23910
rect 22756 23962 22812 23964
rect 22836 23962 22892 23964
rect 22916 23962 22972 23964
rect 22996 23962 23052 23964
rect 22756 23910 22782 23962
rect 22782 23910 22812 23962
rect 22836 23910 22846 23962
rect 22846 23910 22892 23962
rect 22916 23910 22962 23962
rect 22962 23910 22972 23962
rect 22996 23910 23026 23962
rect 23026 23910 23052 23962
rect 22756 23908 22812 23910
rect 22836 23908 22892 23910
rect 22916 23908 22972 23910
rect 22996 23908 23052 23910
rect 3256 23418 3312 23420
rect 3336 23418 3392 23420
rect 3416 23418 3472 23420
rect 3496 23418 3552 23420
rect 3256 23366 3282 23418
rect 3282 23366 3312 23418
rect 3336 23366 3346 23418
rect 3346 23366 3392 23418
rect 3416 23366 3462 23418
rect 3462 23366 3472 23418
rect 3496 23366 3526 23418
rect 3526 23366 3552 23418
rect 3256 23364 3312 23366
rect 3336 23364 3392 23366
rect 3416 23364 3472 23366
rect 3496 23364 3552 23366
rect 6256 23418 6312 23420
rect 6336 23418 6392 23420
rect 6416 23418 6472 23420
rect 6496 23418 6552 23420
rect 6256 23366 6282 23418
rect 6282 23366 6312 23418
rect 6336 23366 6346 23418
rect 6346 23366 6392 23418
rect 6416 23366 6462 23418
rect 6462 23366 6472 23418
rect 6496 23366 6526 23418
rect 6526 23366 6552 23418
rect 6256 23364 6312 23366
rect 6336 23364 6392 23366
rect 6416 23364 6472 23366
rect 6496 23364 6552 23366
rect 9256 23418 9312 23420
rect 9336 23418 9392 23420
rect 9416 23418 9472 23420
rect 9496 23418 9552 23420
rect 9256 23366 9282 23418
rect 9282 23366 9312 23418
rect 9336 23366 9346 23418
rect 9346 23366 9392 23418
rect 9416 23366 9462 23418
rect 9462 23366 9472 23418
rect 9496 23366 9526 23418
rect 9526 23366 9552 23418
rect 9256 23364 9312 23366
rect 9336 23364 9392 23366
rect 9416 23364 9472 23366
rect 9496 23364 9552 23366
rect 12256 23418 12312 23420
rect 12336 23418 12392 23420
rect 12416 23418 12472 23420
rect 12496 23418 12552 23420
rect 12256 23366 12282 23418
rect 12282 23366 12312 23418
rect 12336 23366 12346 23418
rect 12346 23366 12392 23418
rect 12416 23366 12462 23418
rect 12462 23366 12472 23418
rect 12496 23366 12526 23418
rect 12526 23366 12552 23418
rect 12256 23364 12312 23366
rect 12336 23364 12392 23366
rect 12416 23364 12472 23366
rect 12496 23364 12552 23366
rect 15256 23418 15312 23420
rect 15336 23418 15392 23420
rect 15416 23418 15472 23420
rect 15496 23418 15552 23420
rect 15256 23366 15282 23418
rect 15282 23366 15312 23418
rect 15336 23366 15346 23418
rect 15346 23366 15392 23418
rect 15416 23366 15462 23418
rect 15462 23366 15472 23418
rect 15496 23366 15526 23418
rect 15526 23366 15552 23418
rect 15256 23364 15312 23366
rect 15336 23364 15392 23366
rect 15416 23364 15472 23366
rect 15496 23364 15552 23366
rect 18256 23418 18312 23420
rect 18336 23418 18392 23420
rect 18416 23418 18472 23420
rect 18496 23418 18552 23420
rect 18256 23366 18282 23418
rect 18282 23366 18312 23418
rect 18336 23366 18346 23418
rect 18346 23366 18392 23418
rect 18416 23366 18462 23418
rect 18462 23366 18472 23418
rect 18496 23366 18526 23418
rect 18526 23366 18552 23418
rect 18256 23364 18312 23366
rect 18336 23364 18392 23366
rect 18416 23364 18472 23366
rect 18496 23364 18552 23366
rect 21256 23418 21312 23420
rect 21336 23418 21392 23420
rect 21416 23418 21472 23420
rect 21496 23418 21552 23420
rect 21256 23366 21282 23418
rect 21282 23366 21312 23418
rect 21336 23366 21346 23418
rect 21346 23366 21392 23418
rect 21416 23366 21462 23418
rect 21462 23366 21472 23418
rect 21496 23366 21526 23418
rect 21526 23366 21552 23418
rect 21256 23364 21312 23366
rect 21336 23364 21392 23366
rect 21416 23364 21472 23366
rect 21496 23364 21552 23366
rect 1756 22874 1812 22876
rect 1836 22874 1892 22876
rect 1916 22874 1972 22876
rect 1996 22874 2052 22876
rect 1756 22822 1782 22874
rect 1782 22822 1812 22874
rect 1836 22822 1846 22874
rect 1846 22822 1892 22874
rect 1916 22822 1962 22874
rect 1962 22822 1972 22874
rect 1996 22822 2026 22874
rect 2026 22822 2052 22874
rect 1756 22820 1812 22822
rect 1836 22820 1892 22822
rect 1916 22820 1972 22822
rect 1996 22820 2052 22822
rect 4756 22874 4812 22876
rect 4836 22874 4892 22876
rect 4916 22874 4972 22876
rect 4996 22874 5052 22876
rect 4756 22822 4782 22874
rect 4782 22822 4812 22874
rect 4836 22822 4846 22874
rect 4846 22822 4892 22874
rect 4916 22822 4962 22874
rect 4962 22822 4972 22874
rect 4996 22822 5026 22874
rect 5026 22822 5052 22874
rect 4756 22820 4812 22822
rect 4836 22820 4892 22822
rect 4916 22820 4972 22822
rect 4996 22820 5052 22822
rect 7756 22874 7812 22876
rect 7836 22874 7892 22876
rect 7916 22874 7972 22876
rect 7996 22874 8052 22876
rect 7756 22822 7782 22874
rect 7782 22822 7812 22874
rect 7836 22822 7846 22874
rect 7846 22822 7892 22874
rect 7916 22822 7962 22874
rect 7962 22822 7972 22874
rect 7996 22822 8026 22874
rect 8026 22822 8052 22874
rect 7756 22820 7812 22822
rect 7836 22820 7892 22822
rect 7916 22820 7972 22822
rect 7996 22820 8052 22822
rect 10756 22874 10812 22876
rect 10836 22874 10892 22876
rect 10916 22874 10972 22876
rect 10996 22874 11052 22876
rect 10756 22822 10782 22874
rect 10782 22822 10812 22874
rect 10836 22822 10846 22874
rect 10846 22822 10892 22874
rect 10916 22822 10962 22874
rect 10962 22822 10972 22874
rect 10996 22822 11026 22874
rect 11026 22822 11052 22874
rect 10756 22820 10812 22822
rect 10836 22820 10892 22822
rect 10916 22820 10972 22822
rect 10996 22820 11052 22822
rect 13756 22874 13812 22876
rect 13836 22874 13892 22876
rect 13916 22874 13972 22876
rect 13996 22874 14052 22876
rect 13756 22822 13782 22874
rect 13782 22822 13812 22874
rect 13836 22822 13846 22874
rect 13846 22822 13892 22874
rect 13916 22822 13962 22874
rect 13962 22822 13972 22874
rect 13996 22822 14026 22874
rect 14026 22822 14052 22874
rect 13756 22820 13812 22822
rect 13836 22820 13892 22822
rect 13916 22820 13972 22822
rect 13996 22820 14052 22822
rect 16756 22874 16812 22876
rect 16836 22874 16892 22876
rect 16916 22874 16972 22876
rect 16996 22874 17052 22876
rect 16756 22822 16782 22874
rect 16782 22822 16812 22874
rect 16836 22822 16846 22874
rect 16846 22822 16892 22874
rect 16916 22822 16962 22874
rect 16962 22822 16972 22874
rect 16996 22822 17026 22874
rect 17026 22822 17052 22874
rect 16756 22820 16812 22822
rect 16836 22820 16892 22822
rect 16916 22820 16972 22822
rect 16996 22820 17052 22822
rect 19756 22874 19812 22876
rect 19836 22874 19892 22876
rect 19916 22874 19972 22876
rect 19996 22874 20052 22876
rect 19756 22822 19782 22874
rect 19782 22822 19812 22874
rect 19836 22822 19846 22874
rect 19846 22822 19892 22874
rect 19916 22822 19962 22874
rect 19962 22822 19972 22874
rect 19996 22822 20026 22874
rect 20026 22822 20052 22874
rect 19756 22820 19812 22822
rect 19836 22820 19892 22822
rect 19916 22820 19972 22822
rect 19996 22820 20052 22822
rect 22756 22874 22812 22876
rect 22836 22874 22892 22876
rect 22916 22874 22972 22876
rect 22996 22874 23052 22876
rect 22756 22822 22782 22874
rect 22782 22822 22812 22874
rect 22836 22822 22846 22874
rect 22846 22822 22892 22874
rect 22916 22822 22962 22874
rect 22962 22822 22972 22874
rect 22996 22822 23026 22874
rect 23026 22822 23052 22874
rect 22756 22820 22812 22822
rect 22836 22820 22892 22822
rect 22916 22820 22972 22822
rect 22996 22820 23052 22822
rect 3256 22330 3312 22332
rect 3336 22330 3392 22332
rect 3416 22330 3472 22332
rect 3496 22330 3552 22332
rect 3256 22278 3282 22330
rect 3282 22278 3312 22330
rect 3336 22278 3346 22330
rect 3346 22278 3392 22330
rect 3416 22278 3462 22330
rect 3462 22278 3472 22330
rect 3496 22278 3526 22330
rect 3526 22278 3552 22330
rect 3256 22276 3312 22278
rect 3336 22276 3392 22278
rect 3416 22276 3472 22278
rect 3496 22276 3552 22278
rect 6256 22330 6312 22332
rect 6336 22330 6392 22332
rect 6416 22330 6472 22332
rect 6496 22330 6552 22332
rect 6256 22278 6282 22330
rect 6282 22278 6312 22330
rect 6336 22278 6346 22330
rect 6346 22278 6392 22330
rect 6416 22278 6462 22330
rect 6462 22278 6472 22330
rect 6496 22278 6526 22330
rect 6526 22278 6552 22330
rect 6256 22276 6312 22278
rect 6336 22276 6392 22278
rect 6416 22276 6472 22278
rect 6496 22276 6552 22278
rect 9256 22330 9312 22332
rect 9336 22330 9392 22332
rect 9416 22330 9472 22332
rect 9496 22330 9552 22332
rect 9256 22278 9282 22330
rect 9282 22278 9312 22330
rect 9336 22278 9346 22330
rect 9346 22278 9392 22330
rect 9416 22278 9462 22330
rect 9462 22278 9472 22330
rect 9496 22278 9526 22330
rect 9526 22278 9552 22330
rect 9256 22276 9312 22278
rect 9336 22276 9392 22278
rect 9416 22276 9472 22278
rect 9496 22276 9552 22278
rect 12256 22330 12312 22332
rect 12336 22330 12392 22332
rect 12416 22330 12472 22332
rect 12496 22330 12552 22332
rect 12256 22278 12282 22330
rect 12282 22278 12312 22330
rect 12336 22278 12346 22330
rect 12346 22278 12392 22330
rect 12416 22278 12462 22330
rect 12462 22278 12472 22330
rect 12496 22278 12526 22330
rect 12526 22278 12552 22330
rect 12256 22276 12312 22278
rect 12336 22276 12392 22278
rect 12416 22276 12472 22278
rect 12496 22276 12552 22278
rect 15256 22330 15312 22332
rect 15336 22330 15392 22332
rect 15416 22330 15472 22332
rect 15496 22330 15552 22332
rect 15256 22278 15282 22330
rect 15282 22278 15312 22330
rect 15336 22278 15346 22330
rect 15346 22278 15392 22330
rect 15416 22278 15462 22330
rect 15462 22278 15472 22330
rect 15496 22278 15526 22330
rect 15526 22278 15552 22330
rect 15256 22276 15312 22278
rect 15336 22276 15392 22278
rect 15416 22276 15472 22278
rect 15496 22276 15552 22278
rect 18256 22330 18312 22332
rect 18336 22330 18392 22332
rect 18416 22330 18472 22332
rect 18496 22330 18552 22332
rect 18256 22278 18282 22330
rect 18282 22278 18312 22330
rect 18336 22278 18346 22330
rect 18346 22278 18392 22330
rect 18416 22278 18462 22330
rect 18462 22278 18472 22330
rect 18496 22278 18526 22330
rect 18526 22278 18552 22330
rect 18256 22276 18312 22278
rect 18336 22276 18392 22278
rect 18416 22276 18472 22278
rect 18496 22276 18552 22278
rect 21256 22330 21312 22332
rect 21336 22330 21392 22332
rect 21416 22330 21472 22332
rect 21496 22330 21552 22332
rect 21256 22278 21282 22330
rect 21282 22278 21312 22330
rect 21336 22278 21346 22330
rect 21346 22278 21392 22330
rect 21416 22278 21462 22330
rect 21462 22278 21472 22330
rect 21496 22278 21526 22330
rect 21526 22278 21552 22330
rect 21256 22276 21312 22278
rect 21336 22276 21392 22278
rect 21416 22276 21472 22278
rect 21496 22276 21552 22278
rect 1756 21786 1812 21788
rect 1836 21786 1892 21788
rect 1916 21786 1972 21788
rect 1996 21786 2052 21788
rect 1756 21734 1782 21786
rect 1782 21734 1812 21786
rect 1836 21734 1846 21786
rect 1846 21734 1892 21786
rect 1916 21734 1962 21786
rect 1962 21734 1972 21786
rect 1996 21734 2026 21786
rect 2026 21734 2052 21786
rect 1756 21732 1812 21734
rect 1836 21732 1892 21734
rect 1916 21732 1972 21734
rect 1996 21732 2052 21734
rect 4756 21786 4812 21788
rect 4836 21786 4892 21788
rect 4916 21786 4972 21788
rect 4996 21786 5052 21788
rect 4756 21734 4782 21786
rect 4782 21734 4812 21786
rect 4836 21734 4846 21786
rect 4846 21734 4892 21786
rect 4916 21734 4962 21786
rect 4962 21734 4972 21786
rect 4996 21734 5026 21786
rect 5026 21734 5052 21786
rect 4756 21732 4812 21734
rect 4836 21732 4892 21734
rect 4916 21732 4972 21734
rect 4996 21732 5052 21734
rect 7756 21786 7812 21788
rect 7836 21786 7892 21788
rect 7916 21786 7972 21788
rect 7996 21786 8052 21788
rect 7756 21734 7782 21786
rect 7782 21734 7812 21786
rect 7836 21734 7846 21786
rect 7846 21734 7892 21786
rect 7916 21734 7962 21786
rect 7962 21734 7972 21786
rect 7996 21734 8026 21786
rect 8026 21734 8052 21786
rect 7756 21732 7812 21734
rect 7836 21732 7892 21734
rect 7916 21732 7972 21734
rect 7996 21732 8052 21734
rect 10756 21786 10812 21788
rect 10836 21786 10892 21788
rect 10916 21786 10972 21788
rect 10996 21786 11052 21788
rect 10756 21734 10782 21786
rect 10782 21734 10812 21786
rect 10836 21734 10846 21786
rect 10846 21734 10892 21786
rect 10916 21734 10962 21786
rect 10962 21734 10972 21786
rect 10996 21734 11026 21786
rect 11026 21734 11052 21786
rect 10756 21732 10812 21734
rect 10836 21732 10892 21734
rect 10916 21732 10972 21734
rect 10996 21732 11052 21734
rect 13756 21786 13812 21788
rect 13836 21786 13892 21788
rect 13916 21786 13972 21788
rect 13996 21786 14052 21788
rect 13756 21734 13782 21786
rect 13782 21734 13812 21786
rect 13836 21734 13846 21786
rect 13846 21734 13892 21786
rect 13916 21734 13962 21786
rect 13962 21734 13972 21786
rect 13996 21734 14026 21786
rect 14026 21734 14052 21786
rect 13756 21732 13812 21734
rect 13836 21732 13892 21734
rect 13916 21732 13972 21734
rect 13996 21732 14052 21734
rect 16756 21786 16812 21788
rect 16836 21786 16892 21788
rect 16916 21786 16972 21788
rect 16996 21786 17052 21788
rect 16756 21734 16782 21786
rect 16782 21734 16812 21786
rect 16836 21734 16846 21786
rect 16846 21734 16892 21786
rect 16916 21734 16962 21786
rect 16962 21734 16972 21786
rect 16996 21734 17026 21786
rect 17026 21734 17052 21786
rect 16756 21732 16812 21734
rect 16836 21732 16892 21734
rect 16916 21732 16972 21734
rect 16996 21732 17052 21734
rect 19756 21786 19812 21788
rect 19836 21786 19892 21788
rect 19916 21786 19972 21788
rect 19996 21786 20052 21788
rect 19756 21734 19782 21786
rect 19782 21734 19812 21786
rect 19836 21734 19846 21786
rect 19846 21734 19892 21786
rect 19916 21734 19962 21786
rect 19962 21734 19972 21786
rect 19996 21734 20026 21786
rect 20026 21734 20052 21786
rect 19756 21732 19812 21734
rect 19836 21732 19892 21734
rect 19916 21732 19972 21734
rect 19996 21732 20052 21734
rect 22756 21786 22812 21788
rect 22836 21786 22892 21788
rect 22916 21786 22972 21788
rect 22996 21786 23052 21788
rect 22756 21734 22782 21786
rect 22782 21734 22812 21786
rect 22836 21734 22846 21786
rect 22846 21734 22892 21786
rect 22916 21734 22962 21786
rect 22962 21734 22972 21786
rect 22996 21734 23026 21786
rect 23026 21734 23052 21786
rect 22756 21732 22812 21734
rect 22836 21732 22892 21734
rect 22916 21732 22972 21734
rect 22996 21732 23052 21734
rect 3256 21242 3312 21244
rect 3336 21242 3392 21244
rect 3416 21242 3472 21244
rect 3496 21242 3552 21244
rect 3256 21190 3282 21242
rect 3282 21190 3312 21242
rect 3336 21190 3346 21242
rect 3346 21190 3392 21242
rect 3416 21190 3462 21242
rect 3462 21190 3472 21242
rect 3496 21190 3526 21242
rect 3526 21190 3552 21242
rect 3256 21188 3312 21190
rect 3336 21188 3392 21190
rect 3416 21188 3472 21190
rect 3496 21188 3552 21190
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6416 21242 6472 21244
rect 6496 21242 6552 21244
rect 6256 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6416 21190 6462 21242
rect 6462 21190 6472 21242
rect 6496 21190 6526 21242
rect 6526 21190 6552 21242
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 6416 21188 6472 21190
rect 6496 21188 6552 21190
rect 9256 21242 9312 21244
rect 9336 21242 9392 21244
rect 9416 21242 9472 21244
rect 9496 21242 9552 21244
rect 9256 21190 9282 21242
rect 9282 21190 9312 21242
rect 9336 21190 9346 21242
rect 9346 21190 9392 21242
rect 9416 21190 9462 21242
rect 9462 21190 9472 21242
rect 9496 21190 9526 21242
rect 9526 21190 9552 21242
rect 9256 21188 9312 21190
rect 9336 21188 9392 21190
rect 9416 21188 9472 21190
rect 9496 21188 9552 21190
rect 12256 21242 12312 21244
rect 12336 21242 12392 21244
rect 12416 21242 12472 21244
rect 12496 21242 12552 21244
rect 12256 21190 12282 21242
rect 12282 21190 12312 21242
rect 12336 21190 12346 21242
rect 12346 21190 12392 21242
rect 12416 21190 12462 21242
rect 12462 21190 12472 21242
rect 12496 21190 12526 21242
rect 12526 21190 12552 21242
rect 12256 21188 12312 21190
rect 12336 21188 12392 21190
rect 12416 21188 12472 21190
rect 12496 21188 12552 21190
rect 15256 21242 15312 21244
rect 15336 21242 15392 21244
rect 15416 21242 15472 21244
rect 15496 21242 15552 21244
rect 15256 21190 15282 21242
rect 15282 21190 15312 21242
rect 15336 21190 15346 21242
rect 15346 21190 15392 21242
rect 15416 21190 15462 21242
rect 15462 21190 15472 21242
rect 15496 21190 15526 21242
rect 15526 21190 15552 21242
rect 15256 21188 15312 21190
rect 15336 21188 15392 21190
rect 15416 21188 15472 21190
rect 15496 21188 15552 21190
rect 18256 21242 18312 21244
rect 18336 21242 18392 21244
rect 18416 21242 18472 21244
rect 18496 21242 18552 21244
rect 18256 21190 18282 21242
rect 18282 21190 18312 21242
rect 18336 21190 18346 21242
rect 18346 21190 18392 21242
rect 18416 21190 18462 21242
rect 18462 21190 18472 21242
rect 18496 21190 18526 21242
rect 18526 21190 18552 21242
rect 18256 21188 18312 21190
rect 18336 21188 18392 21190
rect 18416 21188 18472 21190
rect 18496 21188 18552 21190
rect 21256 21242 21312 21244
rect 21336 21242 21392 21244
rect 21416 21242 21472 21244
rect 21496 21242 21552 21244
rect 21256 21190 21282 21242
rect 21282 21190 21312 21242
rect 21336 21190 21346 21242
rect 21346 21190 21392 21242
rect 21416 21190 21462 21242
rect 21462 21190 21472 21242
rect 21496 21190 21526 21242
rect 21526 21190 21552 21242
rect 21256 21188 21312 21190
rect 21336 21188 21392 21190
rect 21416 21188 21472 21190
rect 21496 21188 21552 21190
rect 1756 20698 1812 20700
rect 1836 20698 1892 20700
rect 1916 20698 1972 20700
rect 1996 20698 2052 20700
rect 1756 20646 1782 20698
rect 1782 20646 1812 20698
rect 1836 20646 1846 20698
rect 1846 20646 1892 20698
rect 1916 20646 1962 20698
rect 1962 20646 1972 20698
rect 1996 20646 2026 20698
rect 2026 20646 2052 20698
rect 1756 20644 1812 20646
rect 1836 20644 1892 20646
rect 1916 20644 1972 20646
rect 1996 20644 2052 20646
rect 4756 20698 4812 20700
rect 4836 20698 4892 20700
rect 4916 20698 4972 20700
rect 4996 20698 5052 20700
rect 4756 20646 4782 20698
rect 4782 20646 4812 20698
rect 4836 20646 4846 20698
rect 4846 20646 4892 20698
rect 4916 20646 4962 20698
rect 4962 20646 4972 20698
rect 4996 20646 5026 20698
rect 5026 20646 5052 20698
rect 4756 20644 4812 20646
rect 4836 20644 4892 20646
rect 4916 20644 4972 20646
rect 4996 20644 5052 20646
rect 7756 20698 7812 20700
rect 7836 20698 7892 20700
rect 7916 20698 7972 20700
rect 7996 20698 8052 20700
rect 7756 20646 7782 20698
rect 7782 20646 7812 20698
rect 7836 20646 7846 20698
rect 7846 20646 7892 20698
rect 7916 20646 7962 20698
rect 7962 20646 7972 20698
rect 7996 20646 8026 20698
rect 8026 20646 8052 20698
rect 7756 20644 7812 20646
rect 7836 20644 7892 20646
rect 7916 20644 7972 20646
rect 7996 20644 8052 20646
rect 10756 20698 10812 20700
rect 10836 20698 10892 20700
rect 10916 20698 10972 20700
rect 10996 20698 11052 20700
rect 10756 20646 10782 20698
rect 10782 20646 10812 20698
rect 10836 20646 10846 20698
rect 10846 20646 10892 20698
rect 10916 20646 10962 20698
rect 10962 20646 10972 20698
rect 10996 20646 11026 20698
rect 11026 20646 11052 20698
rect 10756 20644 10812 20646
rect 10836 20644 10892 20646
rect 10916 20644 10972 20646
rect 10996 20644 11052 20646
rect 13756 20698 13812 20700
rect 13836 20698 13892 20700
rect 13916 20698 13972 20700
rect 13996 20698 14052 20700
rect 13756 20646 13782 20698
rect 13782 20646 13812 20698
rect 13836 20646 13846 20698
rect 13846 20646 13892 20698
rect 13916 20646 13962 20698
rect 13962 20646 13972 20698
rect 13996 20646 14026 20698
rect 14026 20646 14052 20698
rect 13756 20644 13812 20646
rect 13836 20644 13892 20646
rect 13916 20644 13972 20646
rect 13996 20644 14052 20646
rect 16756 20698 16812 20700
rect 16836 20698 16892 20700
rect 16916 20698 16972 20700
rect 16996 20698 17052 20700
rect 16756 20646 16782 20698
rect 16782 20646 16812 20698
rect 16836 20646 16846 20698
rect 16846 20646 16892 20698
rect 16916 20646 16962 20698
rect 16962 20646 16972 20698
rect 16996 20646 17026 20698
rect 17026 20646 17052 20698
rect 16756 20644 16812 20646
rect 16836 20644 16892 20646
rect 16916 20644 16972 20646
rect 16996 20644 17052 20646
rect 19756 20698 19812 20700
rect 19836 20698 19892 20700
rect 19916 20698 19972 20700
rect 19996 20698 20052 20700
rect 19756 20646 19782 20698
rect 19782 20646 19812 20698
rect 19836 20646 19846 20698
rect 19846 20646 19892 20698
rect 19916 20646 19962 20698
rect 19962 20646 19972 20698
rect 19996 20646 20026 20698
rect 20026 20646 20052 20698
rect 19756 20644 19812 20646
rect 19836 20644 19892 20646
rect 19916 20644 19972 20646
rect 19996 20644 20052 20646
rect 22756 20698 22812 20700
rect 22836 20698 22892 20700
rect 22916 20698 22972 20700
rect 22996 20698 23052 20700
rect 22756 20646 22782 20698
rect 22782 20646 22812 20698
rect 22836 20646 22846 20698
rect 22846 20646 22892 20698
rect 22916 20646 22962 20698
rect 22962 20646 22972 20698
rect 22996 20646 23026 20698
rect 23026 20646 23052 20698
rect 22756 20644 22812 20646
rect 22836 20644 22892 20646
rect 22916 20644 22972 20646
rect 22996 20644 23052 20646
rect 3256 20154 3312 20156
rect 3336 20154 3392 20156
rect 3416 20154 3472 20156
rect 3496 20154 3552 20156
rect 3256 20102 3282 20154
rect 3282 20102 3312 20154
rect 3336 20102 3346 20154
rect 3346 20102 3392 20154
rect 3416 20102 3462 20154
rect 3462 20102 3472 20154
rect 3496 20102 3526 20154
rect 3526 20102 3552 20154
rect 3256 20100 3312 20102
rect 3336 20100 3392 20102
rect 3416 20100 3472 20102
rect 3496 20100 3552 20102
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6416 20154 6472 20156
rect 6496 20154 6552 20156
rect 6256 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6416 20102 6462 20154
rect 6462 20102 6472 20154
rect 6496 20102 6526 20154
rect 6526 20102 6552 20154
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 6416 20100 6472 20102
rect 6496 20100 6552 20102
rect 9256 20154 9312 20156
rect 9336 20154 9392 20156
rect 9416 20154 9472 20156
rect 9496 20154 9552 20156
rect 9256 20102 9282 20154
rect 9282 20102 9312 20154
rect 9336 20102 9346 20154
rect 9346 20102 9392 20154
rect 9416 20102 9462 20154
rect 9462 20102 9472 20154
rect 9496 20102 9526 20154
rect 9526 20102 9552 20154
rect 9256 20100 9312 20102
rect 9336 20100 9392 20102
rect 9416 20100 9472 20102
rect 9496 20100 9552 20102
rect 12256 20154 12312 20156
rect 12336 20154 12392 20156
rect 12416 20154 12472 20156
rect 12496 20154 12552 20156
rect 12256 20102 12282 20154
rect 12282 20102 12312 20154
rect 12336 20102 12346 20154
rect 12346 20102 12392 20154
rect 12416 20102 12462 20154
rect 12462 20102 12472 20154
rect 12496 20102 12526 20154
rect 12526 20102 12552 20154
rect 12256 20100 12312 20102
rect 12336 20100 12392 20102
rect 12416 20100 12472 20102
rect 12496 20100 12552 20102
rect 15256 20154 15312 20156
rect 15336 20154 15392 20156
rect 15416 20154 15472 20156
rect 15496 20154 15552 20156
rect 15256 20102 15282 20154
rect 15282 20102 15312 20154
rect 15336 20102 15346 20154
rect 15346 20102 15392 20154
rect 15416 20102 15462 20154
rect 15462 20102 15472 20154
rect 15496 20102 15526 20154
rect 15526 20102 15552 20154
rect 15256 20100 15312 20102
rect 15336 20100 15392 20102
rect 15416 20100 15472 20102
rect 15496 20100 15552 20102
rect 18256 20154 18312 20156
rect 18336 20154 18392 20156
rect 18416 20154 18472 20156
rect 18496 20154 18552 20156
rect 18256 20102 18282 20154
rect 18282 20102 18312 20154
rect 18336 20102 18346 20154
rect 18346 20102 18392 20154
rect 18416 20102 18462 20154
rect 18462 20102 18472 20154
rect 18496 20102 18526 20154
rect 18526 20102 18552 20154
rect 18256 20100 18312 20102
rect 18336 20100 18392 20102
rect 18416 20100 18472 20102
rect 18496 20100 18552 20102
rect 21256 20154 21312 20156
rect 21336 20154 21392 20156
rect 21416 20154 21472 20156
rect 21496 20154 21552 20156
rect 21256 20102 21282 20154
rect 21282 20102 21312 20154
rect 21336 20102 21346 20154
rect 21346 20102 21392 20154
rect 21416 20102 21462 20154
rect 21462 20102 21472 20154
rect 21496 20102 21526 20154
rect 21526 20102 21552 20154
rect 21256 20100 21312 20102
rect 21336 20100 21392 20102
rect 21416 20100 21472 20102
rect 21496 20100 21552 20102
rect 1756 19610 1812 19612
rect 1836 19610 1892 19612
rect 1916 19610 1972 19612
rect 1996 19610 2052 19612
rect 1756 19558 1782 19610
rect 1782 19558 1812 19610
rect 1836 19558 1846 19610
rect 1846 19558 1892 19610
rect 1916 19558 1962 19610
rect 1962 19558 1972 19610
rect 1996 19558 2026 19610
rect 2026 19558 2052 19610
rect 1756 19556 1812 19558
rect 1836 19556 1892 19558
rect 1916 19556 1972 19558
rect 1996 19556 2052 19558
rect 4756 19610 4812 19612
rect 4836 19610 4892 19612
rect 4916 19610 4972 19612
rect 4996 19610 5052 19612
rect 4756 19558 4782 19610
rect 4782 19558 4812 19610
rect 4836 19558 4846 19610
rect 4846 19558 4892 19610
rect 4916 19558 4962 19610
rect 4962 19558 4972 19610
rect 4996 19558 5026 19610
rect 5026 19558 5052 19610
rect 4756 19556 4812 19558
rect 4836 19556 4892 19558
rect 4916 19556 4972 19558
rect 4996 19556 5052 19558
rect 7756 19610 7812 19612
rect 7836 19610 7892 19612
rect 7916 19610 7972 19612
rect 7996 19610 8052 19612
rect 7756 19558 7782 19610
rect 7782 19558 7812 19610
rect 7836 19558 7846 19610
rect 7846 19558 7892 19610
rect 7916 19558 7962 19610
rect 7962 19558 7972 19610
rect 7996 19558 8026 19610
rect 8026 19558 8052 19610
rect 7756 19556 7812 19558
rect 7836 19556 7892 19558
rect 7916 19556 7972 19558
rect 7996 19556 8052 19558
rect 10756 19610 10812 19612
rect 10836 19610 10892 19612
rect 10916 19610 10972 19612
rect 10996 19610 11052 19612
rect 10756 19558 10782 19610
rect 10782 19558 10812 19610
rect 10836 19558 10846 19610
rect 10846 19558 10892 19610
rect 10916 19558 10962 19610
rect 10962 19558 10972 19610
rect 10996 19558 11026 19610
rect 11026 19558 11052 19610
rect 10756 19556 10812 19558
rect 10836 19556 10892 19558
rect 10916 19556 10972 19558
rect 10996 19556 11052 19558
rect 13756 19610 13812 19612
rect 13836 19610 13892 19612
rect 13916 19610 13972 19612
rect 13996 19610 14052 19612
rect 13756 19558 13782 19610
rect 13782 19558 13812 19610
rect 13836 19558 13846 19610
rect 13846 19558 13892 19610
rect 13916 19558 13962 19610
rect 13962 19558 13972 19610
rect 13996 19558 14026 19610
rect 14026 19558 14052 19610
rect 13756 19556 13812 19558
rect 13836 19556 13892 19558
rect 13916 19556 13972 19558
rect 13996 19556 14052 19558
rect 16756 19610 16812 19612
rect 16836 19610 16892 19612
rect 16916 19610 16972 19612
rect 16996 19610 17052 19612
rect 16756 19558 16782 19610
rect 16782 19558 16812 19610
rect 16836 19558 16846 19610
rect 16846 19558 16892 19610
rect 16916 19558 16962 19610
rect 16962 19558 16972 19610
rect 16996 19558 17026 19610
rect 17026 19558 17052 19610
rect 16756 19556 16812 19558
rect 16836 19556 16892 19558
rect 16916 19556 16972 19558
rect 16996 19556 17052 19558
rect 19756 19610 19812 19612
rect 19836 19610 19892 19612
rect 19916 19610 19972 19612
rect 19996 19610 20052 19612
rect 19756 19558 19782 19610
rect 19782 19558 19812 19610
rect 19836 19558 19846 19610
rect 19846 19558 19892 19610
rect 19916 19558 19962 19610
rect 19962 19558 19972 19610
rect 19996 19558 20026 19610
rect 20026 19558 20052 19610
rect 19756 19556 19812 19558
rect 19836 19556 19892 19558
rect 19916 19556 19972 19558
rect 19996 19556 20052 19558
rect 22756 19610 22812 19612
rect 22836 19610 22892 19612
rect 22916 19610 22972 19612
rect 22996 19610 23052 19612
rect 22756 19558 22782 19610
rect 22782 19558 22812 19610
rect 22836 19558 22846 19610
rect 22846 19558 22892 19610
rect 22916 19558 22962 19610
rect 22962 19558 22972 19610
rect 22996 19558 23026 19610
rect 23026 19558 23052 19610
rect 22756 19556 22812 19558
rect 22836 19556 22892 19558
rect 22916 19556 22972 19558
rect 22996 19556 23052 19558
rect 3256 19066 3312 19068
rect 3336 19066 3392 19068
rect 3416 19066 3472 19068
rect 3496 19066 3552 19068
rect 3256 19014 3282 19066
rect 3282 19014 3312 19066
rect 3336 19014 3346 19066
rect 3346 19014 3392 19066
rect 3416 19014 3462 19066
rect 3462 19014 3472 19066
rect 3496 19014 3526 19066
rect 3526 19014 3552 19066
rect 3256 19012 3312 19014
rect 3336 19012 3392 19014
rect 3416 19012 3472 19014
rect 3496 19012 3552 19014
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6416 19066 6472 19068
rect 6496 19066 6552 19068
rect 6256 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6416 19014 6462 19066
rect 6462 19014 6472 19066
rect 6496 19014 6526 19066
rect 6526 19014 6552 19066
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 6416 19012 6472 19014
rect 6496 19012 6552 19014
rect 9256 19066 9312 19068
rect 9336 19066 9392 19068
rect 9416 19066 9472 19068
rect 9496 19066 9552 19068
rect 9256 19014 9282 19066
rect 9282 19014 9312 19066
rect 9336 19014 9346 19066
rect 9346 19014 9392 19066
rect 9416 19014 9462 19066
rect 9462 19014 9472 19066
rect 9496 19014 9526 19066
rect 9526 19014 9552 19066
rect 9256 19012 9312 19014
rect 9336 19012 9392 19014
rect 9416 19012 9472 19014
rect 9496 19012 9552 19014
rect 12256 19066 12312 19068
rect 12336 19066 12392 19068
rect 12416 19066 12472 19068
rect 12496 19066 12552 19068
rect 12256 19014 12282 19066
rect 12282 19014 12312 19066
rect 12336 19014 12346 19066
rect 12346 19014 12392 19066
rect 12416 19014 12462 19066
rect 12462 19014 12472 19066
rect 12496 19014 12526 19066
rect 12526 19014 12552 19066
rect 12256 19012 12312 19014
rect 12336 19012 12392 19014
rect 12416 19012 12472 19014
rect 12496 19012 12552 19014
rect 15256 19066 15312 19068
rect 15336 19066 15392 19068
rect 15416 19066 15472 19068
rect 15496 19066 15552 19068
rect 15256 19014 15282 19066
rect 15282 19014 15312 19066
rect 15336 19014 15346 19066
rect 15346 19014 15392 19066
rect 15416 19014 15462 19066
rect 15462 19014 15472 19066
rect 15496 19014 15526 19066
rect 15526 19014 15552 19066
rect 15256 19012 15312 19014
rect 15336 19012 15392 19014
rect 15416 19012 15472 19014
rect 15496 19012 15552 19014
rect 18256 19066 18312 19068
rect 18336 19066 18392 19068
rect 18416 19066 18472 19068
rect 18496 19066 18552 19068
rect 18256 19014 18282 19066
rect 18282 19014 18312 19066
rect 18336 19014 18346 19066
rect 18346 19014 18392 19066
rect 18416 19014 18462 19066
rect 18462 19014 18472 19066
rect 18496 19014 18526 19066
rect 18526 19014 18552 19066
rect 18256 19012 18312 19014
rect 18336 19012 18392 19014
rect 18416 19012 18472 19014
rect 18496 19012 18552 19014
rect 21256 19066 21312 19068
rect 21336 19066 21392 19068
rect 21416 19066 21472 19068
rect 21496 19066 21552 19068
rect 21256 19014 21282 19066
rect 21282 19014 21312 19066
rect 21336 19014 21346 19066
rect 21346 19014 21392 19066
rect 21416 19014 21462 19066
rect 21462 19014 21472 19066
rect 21496 19014 21526 19066
rect 21526 19014 21552 19066
rect 21256 19012 21312 19014
rect 21336 19012 21392 19014
rect 21416 19012 21472 19014
rect 21496 19012 21552 19014
rect 1756 18522 1812 18524
rect 1836 18522 1892 18524
rect 1916 18522 1972 18524
rect 1996 18522 2052 18524
rect 1756 18470 1782 18522
rect 1782 18470 1812 18522
rect 1836 18470 1846 18522
rect 1846 18470 1892 18522
rect 1916 18470 1962 18522
rect 1962 18470 1972 18522
rect 1996 18470 2026 18522
rect 2026 18470 2052 18522
rect 1756 18468 1812 18470
rect 1836 18468 1892 18470
rect 1916 18468 1972 18470
rect 1996 18468 2052 18470
rect 4756 18522 4812 18524
rect 4836 18522 4892 18524
rect 4916 18522 4972 18524
rect 4996 18522 5052 18524
rect 4756 18470 4782 18522
rect 4782 18470 4812 18522
rect 4836 18470 4846 18522
rect 4846 18470 4892 18522
rect 4916 18470 4962 18522
rect 4962 18470 4972 18522
rect 4996 18470 5026 18522
rect 5026 18470 5052 18522
rect 4756 18468 4812 18470
rect 4836 18468 4892 18470
rect 4916 18468 4972 18470
rect 4996 18468 5052 18470
rect 7756 18522 7812 18524
rect 7836 18522 7892 18524
rect 7916 18522 7972 18524
rect 7996 18522 8052 18524
rect 7756 18470 7782 18522
rect 7782 18470 7812 18522
rect 7836 18470 7846 18522
rect 7846 18470 7892 18522
rect 7916 18470 7962 18522
rect 7962 18470 7972 18522
rect 7996 18470 8026 18522
rect 8026 18470 8052 18522
rect 7756 18468 7812 18470
rect 7836 18468 7892 18470
rect 7916 18468 7972 18470
rect 7996 18468 8052 18470
rect 10756 18522 10812 18524
rect 10836 18522 10892 18524
rect 10916 18522 10972 18524
rect 10996 18522 11052 18524
rect 10756 18470 10782 18522
rect 10782 18470 10812 18522
rect 10836 18470 10846 18522
rect 10846 18470 10892 18522
rect 10916 18470 10962 18522
rect 10962 18470 10972 18522
rect 10996 18470 11026 18522
rect 11026 18470 11052 18522
rect 10756 18468 10812 18470
rect 10836 18468 10892 18470
rect 10916 18468 10972 18470
rect 10996 18468 11052 18470
rect 13756 18522 13812 18524
rect 13836 18522 13892 18524
rect 13916 18522 13972 18524
rect 13996 18522 14052 18524
rect 13756 18470 13782 18522
rect 13782 18470 13812 18522
rect 13836 18470 13846 18522
rect 13846 18470 13892 18522
rect 13916 18470 13962 18522
rect 13962 18470 13972 18522
rect 13996 18470 14026 18522
rect 14026 18470 14052 18522
rect 13756 18468 13812 18470
rect 13836 18468 13892 18470
rect 13916 18468 13972 18470
rect 13996 18468 14052 18470
rect 16756 18522 16812 18524
rect 16836 18522 16892 18524
rect 16916 18522 16972 18524
rect 16996 18522 17052 18524
rect 16756 18470 16782 18522
rect 16782 18470 16812 18522
rect 16836 18470 16846 18522
rect 16846 18470 16892 18522
rect 16916 18470 16962 18522
rect 16962 18470 16972 18522
rect 16996 18470 17026 18522
rect 17026 18470 17052 18522
rect 16756 18468 16812 18470
rect 16836 18468 16892 18470
rect 16916 18468 16972 18470
rect 16996 18468 17052 18470
rect 19756 18522 19812 18524
rect 19836 18522 19892 18524
rect 19916 18522 19972 18524
rect 19996 18522 20052 18524
rect 19756 18470 19782 18522
rect 19782 18470 19812 18522
rect 19836 18470 19846 18522
rect 19846 18470 19892 18522
rect 19916 18470 19962 18522
rect 19962 18470 19972 18522
rect 19996 18470 20026 18522
rect 20026 18470 20052 18522
rect 19756 18468 19812 18470
rect 19836 18468 19892 18470
rect 19916 18468 19972 18470
rect 19996 18468 20052 18470
rect 22756 18522 22812 18524
rect 22836 18522 22892 18524
rect 22916 18522 22972 18524
rect 22996 18522 23052 18524
rect 22756 18470 22782 18522
rect 22782 18470 22812 18522
rect 22836 18470 22846 18522
rect 22846 18470 22892 18522
rect 22916 18470 22962 18522
rect 22962 18470 22972 18522
rect 22996 18470 23026 18522
rect 23026 18470 23052 18522
rect 22756 18468 22812 18470
rect 22836 18468 22892 18470
rect 22916 18468 22972 18470
rect 22996 18468 23052 18470
rect 3256 17978 3312 17980
rect 3336 17978 3392 17980
rect 3416 17978 3472 17980
rect 3496 17978 3552 17980
rect 3256 17926 3282 17978
rect 3282 17926 3312 17978
rect 3336 17926 3346 17978
rect 3346 17926 3392 17978
rect 3416 17926 3462 17978
rect 3462 17926 3472 17978
rect 3496 17926 3526 17978
rect 3526 17926 3552 17978
rect 3256 17924 3312 17926
rect 3336 17924 3392 17926
rect 3416 17924 3472 17926
rect 3496 17924 3552 17926
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6416 17978 6472 17980
rect 6496 17978 6552 17980
rect 6256 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6416 17926 6462 17978
rect 6462 17926 6472 17978
rect 6496 17926 6526 17978
rect 6526 17926 6552 17978
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 6416 17924 6472 17926
rect 6496 17924 6552 17926
rect 9256 17978 9312 17980
rect 9336 17978 9392 17980
rect 9416 17978 9472 17980
rect 9496 17978 9552 17980
rect 9256 17926 9282 17978
rect 9282 17926 9312 17978
rect 9336 17926 9346 17978
rect 9346 17926 9392 17978
rect 9416 17926 9462 17978
rect 9462 17926 9472 17978
rect 9496 17926 9526 17978
rect 9526 17926 9552 17978
rect 9256 17924 9312 17926
rect 9336 17924 9392 17926
rect 9416 17924 9472 17926
rect 9496 17924 9552 17926
rect 12256 17978 12312 17980
rect 12336 17978 12392 17980
rect 12416 17978 12472 17980
rect 12496 17978 12552 17980
rect 12256 17926 12282 17978
rect 12282 17926 12312 17978
rect 12336 17926 12346 17978
rect 12346 17926 12392 17978
rect 12416 17926 12462 17978
rect 12462 17926 12472 17978
rect 12496 17926 12526 17978
rect 12526 17926 12552 17978
rect 12256 17924 12312 17926
rect 12336 17924 12392 17926
rect 12416 17924 12472 17926
rect 12496 17924 12552 17926
rect 15256 17978 15312 17980
rect 15336 17978 15392 17980
rect 15416 17978 15472 17980
rect 15496 17978 15552 17980
rect 15256 17926 15282 17978
rect 15282 17926 15312 17978
rect 15336 17926 15346 17978
rect 15346 17926 15392 17978
rect 15416 17926 15462 17978
rect 15462 17926 15472 17978
rect 15496 17926 15526 17978
rect 15526 17926 15552 17978
rect 15256 17924 15312 17926
rect 15336 17924 15392 17926
rect 15416 17924 15472 17926
rect 15496 17924 15552 17926
rect 18256 17978 18312 17980
rect 18336 17978 18392 17980
rect 18416 17978 18472 17980
rect 18496 17978 18552 17980
rect 18256 17926 18282 17978
rect 18282 17926 18312 17978
rect 18336 17926 18346 17978
rect 18346 17926 18392 17978
rect 18416 17926 18462 17978
rect 18462 17926 18472 17978
rect 18496 17926 18526 17978
rect 18526 17926 18552 17978
rect 18256 17924 18312 17926
rect 18336 17924 18392 17926
rect 18416 17924 18472 17926
rect 18496 17924 18552 17926
rect 21256 17978 21312 17980
rect 21336 17978 21392 17980
rect 21416 17978 21472 17980
rect 21496 17978 21552 17980
rect 21256 17926 21282 17978
rect 21282 17926 21312 17978
rect 21336 17926 21346 17978
rect 21346 17926 21392 17978
rect 21416 17926 21462 17978
rect 21462 17926 21472 17978
rect 21496 17926 21526 17978
rect 21526 17926 21552 17978
rect 21256 17924 21312 17926
rect 21336 17924 21392 17926
rect 21416 17924 21472 17926
rect 21496 17924 21552 17926
rect 1756 17434 1812 17436
rect 1836 17434 1892 17436
rect 1916 17434 1972 17436
rect 1996 17434 2052 17436
rect 1756 17382 1782 17434
rect 1782 17382 1812 17434
rect 1836 17382 1846 17434
rect 1846 17382 1892 17434
rect 1916 17382 1962 17434
rect 1962 17382 1972 17434
rect 1996 17382 2026 17434
rect 2026 17382 2052 17434
rect 1756 17380 1812 17382
rect 1836 17380 1892 17382
rect 1916 17380 1972 17382
rect 1996 17380 2052 17382
rect 4756 17434 4812 17436
rect 4836 17434 4892 17436
rect 4916 17434 4972 17436
rect 4996 17434 5052 17436
rect 4756 17382 4782 17434
rect 4782 17382 4812 17434
rect 4836 17382 4846 17434
rect 4846 17382 4892 17434
rect 4916 17382 4962 17434
rect 4962 17382 4972 17434
rect 4996 17382 5026 17434
rect 5026 17382 5052 17434
rect 4756 17380 4812 17382
rect 4836 17380 4892 17382
rect 4916 17380 4972 17382
rect 4996 17380 5052 17382
rect 7756 17434 7812 17436
rect 7836 17434 7892 17436
rect 7916 17434 7972 17436
rect 7996 17434 8052 17436
rect 7756 17382 7782 17434
rect 7782 17382 7812 17434
rect 7836 17382 7846 17434
rect 7846 17382 7892 17434
rect 7916 17382 7962 17434
rect 7962 17382 7972 17434
rect 7996 17382 8026 17434
rect 8026 17382 8052 17434
rect 7756 17380 7812 17382
rect 7836 17380 7892 17382
rect 7916 17380 7972 17382
rect 7996 17380 8052 17382
rect 10756 17434 10812 17436
rect 10836 17434 10892 17436
rect 10916 17434 10972 17436
rect 10996 17434 11052 17436
rect 10756 17382 10782 17434
rect 10782 17382 10812 17434
rect 10836 17382 10846 17434
rect 10846 17382 10892 17434
rect 10916 17382 10962 17434
rect 10962 17382 10972 17434
rect 10996 17382 11026 17434
rect 11026 17382 11052 17434
rect 10756 17380 10812 17382
rect 10836 17380 10892 17382
rect 10916 17380 10972 17382
rect 10996 17380 11052 17382
rect 13756 17434 13812 17436
rect 13836 17434 13892 17436
rect 13916 17434 13972 17436
rect 13996 17434 14052 17436
rect 13756 17382 13782 17434
rect 13782 17382 13812 17434
rect 13836 17382 13846 17434
rect 13846 17382 13892 17434
rect 13916 17382 13962 17434
rect 13962 17382 13972 17434
rect 13996 17382 14026 17434
rect 14026 17382 14052 17434
rect 13756 17380 13812 17382
rect 13836 17380 13892 17382
rect 13916 17380 13972 17382
rect 13996 17380 14052 17382
rect 16756 17434 16812 17436
rect 16836 17434 16892 17436
rect 16916 17434 16972 17436
rect 16996 17434 17052 17436
rect 16756 17382 16782 17434
rect 16782 17382 16812 17434
rect 16836 17382 16846 17434
rect 16846 17382 16892 17434
rect 16916 17382 16962 17434
rect 16962 17382 16972 17434
rect 16996 17382 17026 17434
rect 17026 17382 17052 17434
rect 16756 17380 16812 17382
rect 16836 17380 16892 17382
rect 16916 17380 16972 17382
rect 16996 17380 17052 17382
rect 19756 17434 19812 17436
rect 19836 17434 19892 17436
rect 19916 17434 19972 17436
rect 19996 17434 20052 17436
rect 19756 17382 19782 17434
rect 19782 17382 19812 17434
rect 19836 17382 19846 17434
rect 19846 17382 19892 17434
rect 19916 17382 19962 17434
rect 19962 17382 19972 17434
rect 19996 17382 20026 17434
rect 20026 17382 20052 17434
rect 19756 17380 19812 17382
rect 19836 17380 19892 17382
rect 19916 17380 19972 17382
rect 19996 17380 20052 17382
rect 22756 17434 22812 17436
rect 22836 17434 22892 17436
rect 22916 17434 22972 17436
rect 22996 17434 23052 17436
rect 22756 17382 22782 17434
rect 22782 17382 22812 17434
rect 22836 17382 22846 17434
rect 22846 17382 22892 17434
rect 22916 17382 22962 17434
rect 22962 17382 22972 17434
rect 22996 17382 23026 17434
rect 23026 17382 23052 17434
rect 22756 17380 22812 17382
rect 22836 17380 22892 17382
rect 22916 17380 22972 17382
rect 22996 17380 23052 17382
rect 3256 16890 3312 16892
rect 3336 16890 3392 16892
rect 3416 16890 3472 16892
rect 3496 16890 3552 16892
rect 3256 16838 3282 16890
rect 3282 16838 3312 16890
rect 3336 16838 3346 16890
rect 3346 16838 3392 16890
rect 3416 16838 3462 16890
rect 3462 16838 3472 16890
rect 3496 16838 3526 16890
rect 3526 16838 3552 16890
rect 3256 16836 3312 16838
rect 3336 16836 3392 16838
rect 3416 16836 3472 16838
rect 3496 16836 3552 16838
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6416 16890 6472 16892
rect 6496 16890 6552 16892
rect 6256 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6416 16838 6462 16890
rect 6462 16838 6472 16890
rect 6496 16838 6526 16890
rect 6526 16838 6552 16890
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6416 16836 6472 16838
rect 6496 16836 6552 16838
rect 9256 16890 9312 16892
rect 9336 16890 9392 16892
rect 9416 16890 9472 16892
rect 9496 16890 9552 16892
rect 9256 16838 9282 16890
rect 9282 16838 9312 16890
rect 9336 16838 9346 16890
rect 9346 16838 9392 16890
rect 9416 16838 9462 16890
rect 9462 16838 9472 16890
rect 9496 16838 9526 16890
rect 9526 16838 9552 16890
rect 9256 16836 9312 16838
rect 9336 16836 9392 16838
rect 9416 16836 9472 16838
rect 9496 16836 9552 16838
rect 12256 16890 12312 16892
rect 12336 16890 12392 16892
rect 12416 16890 12472 16892
rect 12496 16890 12552 16892
rect 12256 16838 12282 16890
rect 12282 16838 12312 16890
rect 12336 16838 12346 16890
rect 12346 16838 12392 16890
rect 12416 16838 12462 16890
rect 12462 16838 12472 16890
rect 12496 16838 12526 16890
rect 12526 16838 12552 16890
rect 12256 16836 12312 16838
rect 12336 16836 12392 16838
rect 12416 16836 12472 16838
rect 12496 16836 12552 16838
rect 15256 16890 15312 16892
rect 15336 16890 15392 16892
rect 15416 16890 15472 16892
rect 15496 16890 15552 16892
rect 15256 16838 15282 16890
rect 15282 16838 15312 16890
rect 15336 16838 15346 16890
rect 15346 16838 15392 16890
rect 15416 16838 15462 16890
rect 15462 16838 15472 16890
rect 15496 16838 15526 16890
rect 15526 16838 15552 16890
rect 15256 16836 15312 16838
rect 15336 16836 15392 16838
rect 15416 16836 15472 16838
rect 15496 16836 15552 16838
rect 18256 16890 18312 16892
rect 18336 16890 18392 16892
rect 18416 16890 18472 16892
rect 18496 16890 18552 16892
rect 18256 16838 18282 16890
rect 18282 16838 18312 16890
rect 18336 16838 18346 16890
rect 18346 16838 18392 16890
rect 18416 16838 18462 16890
rect 18462 16838 18472 16890
rect 18496 16838 18526 16890
rect 18526 16838 18552 16890
rect 18256 16836 18312 16838
rect 18336 16836 18392 16838
rect 18416 16836 18472 16838
rect 18496 16836 18552 16838
rect 21256 16890 21312 16892
rect 21336 16890 21392 16892
rect 21416 16890 21472 16892
rect 21496 16890 21552 16892
rect 21256 16838 21282 16890
rect 21282 16838 21312 16890
rect 21336 16838 21346 16890
rect 21346 16838 21392 16890
rect 21416 16838 21462 16890
rect 21462 16838 21472 16890
rect 21496 16838 21526 16890
rect 21526 16838 21552 16890
rect 21256 16836 21312 16838
rect 21336 16836 21392 16838
rect 21416 16836 21472 16838
rect 21496 16836 21552 16838
rect 1756 16346 1812 16348
rect 1836 16346 1892 16348
rect 1916 16346 1972 16348
rect 1996 16346 2052 16348
rect 1756 16294 1782 16346
rect 1782 16294 1812 16346
rect 1836 16294 1846 16346
rect 1846 16294 1892 16346
rect 1916 16294 1962 16346
rect 1962 16294 1972 16346
rect 1996 16294 2026 16346
rect 2026 16294 2052 16346
rect 1756 16292 1812 16294
rect 1836 16292 1892 16294
rect 1916 16292 1972 16294
rect 1996 16292 2052 16294
rect 4756 16346 4812 16348
rect 4836 16346 4892 16348
rect 4916 16346 4972 16348
rect 4996 16346 5052 16348
rect 4756 16294 4782 16346
rect 4782 16294 4812 16346
rect 4836 16294 4846 16346
rect 4846 16294 4892 16346
rect 4916 16294 4962 16346
rect 4962 16294 4972 16346
rect 4996 16294 5026 16346
rect 5026 16294 5052 16346
rect 4756 16292 4812 16294
rect 4836 16292 4892 16294
rect 4916 16292 4972 16294
rect 4996 16292 5052 16294
rect 7756 16346 7812 16348
rect 7836 16346 7892 16348
rect 7916 16346 7972 16348
rect 7996 16346 8052 16348
rect 7756 16294 7782 16346
rect 7782 16294 7812 16346
rect 7836 16294 7846 16346
rect 7846 16294 7892 16346
rect 7916 16294 7962 16346
rect 7962 16294 7972 16346
rect 7996 16294 8026 16346
rect 8026 16294 8052 16346
rect 7756 16292 7812 16294
rect 7836 16292 7892 16294
rect 7916 16292 7972 16294
rect 7996 16292 8052 16294
rect 10756 16346 10812 16348
rect 10836 16346 10892 16348
rect 10916 16346 10972 16348
rect 10996 16346 11052 16348
rect 10756 16294 10782 16346
rect 10782 16294 10812 16346
rect 10836 16294 10846 16346
rect 10846 16294 10892 16346
rect 10916 16294 10962 16346
rect 10962 16294 10972 16346
rect 10996 16294 11026 16346
rect 11026 16294 11052 16346
rect 10756 16292 10812 16294
rect 10836 16292 10892 16294
rect 10916 16292 10972 16294
rect 10996 16292 11052 16294
rect 13756 16346 13812 16348
rect 13836 16346 13892 16348
rect 13916 16346 13972 16348
rect 13996 16346 14052 16348
rect 13756 16294 13782 16346
rect 13782 16294 13812 16346
rect 13836 16294 13846 16346
rect 13846 16294 13892 16346
rect 13916 16294 13962 16346
rect 13962 16294 13972 16346
rect 13996 16294 14026 16346
rect 14026 16294 14052 16346
rect 13756 16292 13812 16294
rect 13836 16292 13892 16294
rect 13916 16292 13972 16294
rect 13996 16292 14052 16294
rect 3256 15802 3312 15804
rect 3336 15802 3392 15804
rect 3416 15802 3472 15804
rect 3496 15802 3552 15804
rect 3256 15750 3282 15802
rect 3282 15750 3312 15802
rect 3336 15750 3346 15802
rect 3346 15750 3392 15802
rect 3416 15750 3462 15802
rect 3462 15750 3472 15802
rect 3496 15750 3526 15802
rect 3526 15750 3552 15802
rect 3256 15748 3312 15750
rect 3336 15748 3392 15750
rect 3416 15748 3472 15750
rect 3496 15748 3552 15750
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6416 15802 6472 15804
rect 6496 15802 6552 15804
rect 6256 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6416 15750 6462 15802
rect 6462 15750 6472 15802
rect 6496 15750 6526 15802
rect 6526 15750 6552 15802
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6416 15748 6472 15750
rect 6496 15748 6552 15750
rect 9256 15802 9312 15804
rect 9336 15802 9392 15804
rect 9416 15802 9472 15804
rect 9496 15802 9552 15804
rect 9256 15750 9282 15802
rect 9282 15750 9312 15802
rect 9336 15750 9346 15802
rect 9346 15750 9392 15802
rect 9416 15750 9462 15802
rect 9462 15750 9472 15802
rect 9496 15750 9526 15802
rect 9526 15750 9552 15802
rect 9256 15748 9312 15750
rect 9336 15748 9392 15750
rect 9416 15748 9472 15750
rect 9496 15748 9552 15750
rect 12256 15802 12312 15804
rect 12336 15802 12392 15804
rect 12416 15802 12472 15804
rect 12496 15802 12552 15804
rect 12256 15750 12282 15802
rect 12282 15750 12312 15802
rect 12336 15750 12346 15802
rect 12346 15750 12392 15802
rect 12416 15750 12462 15802
rect 12462 15750 12472 15802
rect 12496 15750 12526 15802
rect 12526 15750 12552 15802
rect 12256 15748 12312 15750
rect 12336 15748 12392 15750
rect 12416 15748 12472 15750
rect 12496 15748 12552 15750
rect 1756 15258 1812 15260
rect 1836 15258 1892 15260
rect 1916 15258 1972 15260
rect 1996 15258 2052 15260
rect 1756 15206 1782 15258
rect 1782 15206 1812 15258
rect 1836 15206 1846 15258
rect 1846 15206 1892 15258
rect 1916 15206 1962 15258
rect 1962 15206 1972 15258
rect 1996 15206 2026 15258
rect 2026 15206 2052 15258
rect 1756 15204 1812 15206
rect 1836 15204 1892 15206
rect 1916 15204 1972 15206
rect 1996 15204 2052 15206
rect 4756 15258 4812 15260
rect 4836 15258 4892 15260
rect 4916 15258 4972 15260
rect 4996 15258 5052 15260
rect 4756 15206 4782 15258
rect 4782 15206 4812 15258
rect 4836 15206 4846 15258
rect 4846 15206 4892 15258
rect 4916 15206 4962 15258
rect 4962 15206 4972 15258
rect 4996 15206 5026 15258
rect 5026 15206 5052 15258
rect 4756 15204 4812 15206
rect 4836 15204 4892 15206
rect 4916 15204 4972 15206
rect 4996 15204 5052 15206
rect 7756 15258 7812 15260
rect 7836 15258 7892 15260
rect 7916 15258 7972 15260
rect 7996 15258 8052 15260
rect 7756 15206 7782 15258
rect 7782 15206 7812 15258
rect 7836 15206 7846 15258
rect 7846 15206 7892 15258
rect 7916 15206 7962 15258
rect 7962 15206 7972 15258
rect 7996 15206 8026 15258
rect 8026 15206 8052 15258
rect 7756 15204 7812 15206
rect 7836 15204 7892 15206
rect 7916 15204 7972 15206
rect 7996 15204 8052 15206
rect 10756 15258 10812 15260
rect 10836 15258 10892 15260
rect 10916 15258 10972 15260
rect 10996 15258 11052 15260
rect 10756 15206 10782 15258
rect 10782 15206 10812 15258
rect 10836 15206 10846 15258
rect 10846 15206 10892 15258
rect 10916 15206 10962 15258
rect 10962 15206 10972 15258
rect 10996 15206 11026 15258
rect 11026 15206 11052 15258
rect 10756 15204 10812 15206
rect 10836 15204 10892 15206
rect 10916 15204 10972 15206
rect 10996 15204 11052 15206
rect 3256 14714 3312 14716
rect 3336 14714 3392 14716
rect 3416 14714 3472 14716
rect 3496 14714 3552 14716
rect 3256 14662 3282 14714
rect 3282 14662 3312 14714
rect 3336 14662 3346 14714
rect 3346 14662 3392 14714
rect 3416 14662 3462 14714
rect 3462 14662 3472 14714
rect 3496 14662 3526 14714
rect 3526 14662 3552 14714
rect 3256 14660 3312 14662
rect 3336 14660 3392 14662
rect 3416 14660 3472 14662
rect 3496 14660 3552 14662
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6416 14714 6472 14716
rect 6496 14714 6552 14716
rect 6256 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6416 14662 6462 14714
rect 6462 14662 6472 14714
rect 6496 14662 6526 14714
rect 6526 14662 6552 14714
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6416 14660 6472 14662
rect 6496 14660 6552 14662
rect 9256 14714 9312 14716
rect 9336 14714 9392 14716
rect 9416 14714 9472 14716
rect 9496 14714 9552 14716
rect 9256 14662 9282 14714
rect 9282 14662 9312 14714
rect 9336 14662 9346 14714
rect 9346 14662 9392 14714
rect 9416 14662 9462 14714
rect 9462 14662 9472 14714
rect 9496 14662 9526 14714
rect 9526 14662 9552 14714
rect 9256 14660 9312 14662
rect 9336 14660 9392 14662
rect 9416 14660 9472 14662
rect 9496 14660 9552 14662
rect 12256 14714 12312 14716
rect 12336 14714 12392 14716
rect 12416 14714 12472 14716
rect 12496 14714 12552 14716
rect 12256 14662 12282 14714
rect 12282 14662 12312 14714
rect 12336 14662 12346 14714
rect 12346 14662 12392 14714
rect 12416 14662 12462 14714
rect 12462 14662 12472 14714
rect 12496 14662 12526 14714
rect 12526 14662 12552 14714
rect 12256 14660 12312 14662
rect 12336 14660 12392 14662
rect 12416 14660 12472 14662
rect 12496 14660 12552 14662
rect 1756 14170 1812 14172
rect 1836 14170 1892 14172
rect 1916 14170 1972 14172
rect 1996 14170 2052 14172
rect 1756 14118 1782 14170
rect 1782 14118 1812 14170
rect 1836 14118 1846 14170
rect 1846 14118 1892 14170
rect 1916 14118 1962 14170
rect 1962 14118 1972 14170
rect 1996 14118 2026 14170
rect 2026 14118 2052 14170
rect 1756 14116 1812 14118
rect 1836 14116 1892 14118
rect 1916 14116 1972 14118
rect 1996 14116 2052 14118
rect 4756 14170 4812 14172
rect 4836 14170 4892 14172
rect 4916 14170 4972 14172
rect 4996 14170 5052 14172
rect 4756 14118 4782 14170
rect 4782 14118 4812 14170
rect 4836 14118 4846 14170
rect 4846 14118 4892 14170
rect 4916 14118 4962 14170
rect 4962 14118 4972 14170
rect 4996 14118 5026 14170
rect 5026 14118 5052 14170
rect 4756 14116 4812 14118
rect 4836 14116 4892 14118
rect 4916 14116 4972 14118
rect 4996 14116 5052 14118
rect 7756 14170 7812 14172
rect 7836 14170 7892 14172
rect 7916 14170 7972 14172
rect 7996 14170 8052 14172
rect 7756 14118 7782 14170
rect 7782 14118 7812 14170
rect 7836 14118 7846 14170
rect 7846 14118 7892 14170
rect 7916 14118 7962 14170
rect 7962 14118 7972 14170
rect 7996 14118 8026 14170
rect 8026 14118 8052 14170
rect 7756 14116 7812 14118
rect 7836 14116 7892 14118
rect 7916 14116 7972 14118
rect 7996 14116 8052 14118
rect 10756 14170 10812 14172
rect 10836 14170 10892 14172
rect 10916 14170 10972 14172
rect 10996 14170 11052 14172
rect 10756 14118 10782 14170
rect 10782 14118 10812 14170
rect 10836 14118 10846 14170
rect 10846 14118 10892 14170
rect 10916 14118 10962 14170
rect 10962 14118 10972 14170
rect 10996 14118 11026 14170
rect 11026 14118 11052 14170
rect 10756 14116 10812 14118
rect 10836 14116 10892 14118
rect 10916 14116 10972 14118
rect 10996 14116 11052 14118
rect 8482 13932 8538 13968
rect 8482 13912 8484 13932
rect 8484 13912 8536 13932
rect 8536 13912 8538 13932
rect 110 13640 166 13696
rect 3256 13626 3312 13628
rect 3336 13626 3392 13628
rect 3416 13626 3472 13628
rect 3496 13626 3552 13628
rect 3256 13574 3282 13626
rect 3282 13574 3312 13626
rect 3336 13574 3346 13626
rect 3346 13574 3392 13626
rect 3416 13574 3462 13626
rect 3462 13574 3472 13626
rect 3496 13574 3526 13626
rect 3526 13574 3552 13626
rect 3256 13572 3312 13574
rect 3336 13572 3392 13574
rect 3416 13572 3472 13574
rect 3496 13572 3552 13574
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6416 13626 6472 13628
rect 6496 13626 6552 13628
rect 6256 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6416 13574 6462 13626
rect 6462 13574 6472 13626
rect 6496 13574 6526 13626
rect 6526 13574 6552 13626
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6416 13572 6472 13574
rect 6496 13572 6552 13574
rect 1756 13082 1812 13084
rect 1836 13082 1892 13084
rect 1916 13082 1972 13084
rect 1996 13082 2052 13084
rect 1756 13030 1782 13082
rect 1782 13030 1812 13082
rect 1836 13030 1846 13082
rect 1846 13030 1892 13082
rect 1916 13030 1962 13082
rect 1962 13030 1972 13082
rect 1996 13030 2026 13082
rect 2026 13030 2052 13082
rect 1756 13028 1812 13030
rect 1836 13028 1892 13030
rect 1916 13028 1972 13030
rect 1996 13028 2052 13030
rect 4756 13082 4812 13084
rect 4836 13082 4892 13084
rect 4916 13082 4972 13084
rect 4996 13082 5052 13084
rect 4756 13030 4782 13082
rect 4782 13030 4812 13082
rect 4836 13030 4846 13082
rect 4846 13030 4892 13082
rect 4916 13030 4962 13082
rect 4962 13030 4972 13082
rect 4996 13030 5026 13082
rect 5026 13030 5052 13082
rect 4756 13028 4812 13030
rect 4836 13028 4892 13030
rect 4916 13028 4972 13030
rect 4996 13028 5052 13030
rect 7756 13082 7812 13084
rect 7836 13082 7892 13084
rect 7916 13082 7972 13084
rect 7996 13082 8052 13084
rect 7756 13030 7782 13082
rect 7782 13030 7812 13082
rect 7836 13030 7846 13082
rect 7846 13030 7892 13082
rect 7916 13030 7962 13082
rect 7962 13030 7972 13082
rect 7996 13030 8026 13082
rect 8026 13030 8052 13082
rect 7756 13028 7812 13030
rect 7836 13028 7892 13030
rect 7916 13028 7972 13030
rect 7996 13028 8052 13030
rect 110 12688 166 12744
rect 3256 12538 3312 12540
rect 3336 12538 3392 12540
rect 3416 12538 3472 12540
rect 3496 12538 3552 12540
rect 3256 12486 3282 12538
rect 3282 12486 3312 12538
rect 3336 12486 3346 12538
rect 3346 12486 3392 12538
rect 3416 12486 3462 12538
rect 3462 12486 3472 12538
rect 3496 12486 3526 12538
rect 3526 12486 3552 12538
rect 3256 12484 3312 12486
rect 3336 12484 3392 12486
rect 3416 12484 3472 12486
rect 3496 12484 3552 12486
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6416 12538 6472 12540
rect 6496 12538 6552 12540
rect 6256 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6416 12486 6462 12538
rect 6462 12486 6472 12538
rect 6496 12486 6526 12538
rect 6526 12486 6552 12538
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6416 12484 6472 12486
rect 6496 12484 6552 12486
rect 1756 11994 1812 11996
rect 1836 11994 1892 11996
rect 1916 11994 1972 11996
rect 1996 11994 2052 11996
rect 1756 11942 1782 11994
rect 1782 11942 1812 11994
rect 1836 11942 1846 11994
rect 1846 11942 1892 11994
rect 1916 11942 1962 11994
rect 1962 11942 1972 11994
rect 1996 11942 2026 11994
rect 2026 11942 2052 11994
rect 1756 11940 1812 11942
rect 1836 11940 1892 11942
rect 1916 11940 1972 11942
rect 1996 11940 2052 11942
rect 4756 11994 4812 11996
rect 4836 11994 4892 11996
rect 4916 11994 4972 11996
rect 4996 11994 5052 11996
rect 4756 11942 4782 11994
rect 4782 11942 4812 11994
rect 4836 11942 4846 11994
rect 4846 11942 4892 11994
rect 4916 11942 4962 11994
rect 4962 11942 4972 11994
rect 4996 11942 5026 11994
rect 5026 11942 5052 11994
rect 4756 11940 4812 11942
rect 4836 11940 4892 11942
rect 4916 11940 4972 11942
rect 4996 11940 5052 11942
rect 7756 11994 7812 11996
rect 7836 11994 7892 11996
rect 7916 11994 7972 11996
rect 7996 11994 8052 11996
rect 7756 11942 7782 11994
rect 7782 11942 7812 11994
rect 7836 11942 7846 11994
rect 7846 11942 7892 11994
rect 7916 11942 7962 11994
rect 7962 11942 7972 11994
rect 7996 11942 8026 11994
rect 8026 11942 8052 11994
rect 7756 11940 7812 11942
rect 7836 11940 7892 11942
rect 7916 11940 7972 11942
rect 7996 11940 8052 11942
rect 3256 11450 3312 11452
rect 3336 11450 3392 11452
rect 3416 11450 3472 11452
rect 3496 11450 3552 11452
rect 3256 11398 3282 11450
rect 3282 11398 3312 11450
rect 3336 11398 3346 11450
rect 3346 11398 3392 11450
rect 3416 11398 3462 11450
rect 3462 11398 3472 11450
rect 3496 11398 3526 11450
rect 3526 11398 3552 11450
rect 3256 11396 3312 11398
rect 3336 11396 3392 11398
rect 3416 11396 3472 11398
rect 3496 11396 3552 11398
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6416 11450 6472 11452
rect 6496 11450 6552 11452
rect 6256 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6416 11398 6462 11450
rect 6462 11398 6472 11450
rect 6496 11398 6526 11450
rect 6526 11398 6552 11450
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6416 11396 6472 11398
rect 6496 11396 6552 11398
rect 1756 10906 1812 10908
rect 1836 10906 1892 10908
rect 1916 10906 1972 10908
rect 1996 10906 2052 10908
rect 1756 10854 1782 10906
rect 1782 10854 1812 10906
rect 1836 10854 1846 10906
rect 1846 10854 1892 10906
rect 1916 10854 1962 10906
rect 1962 10854 1972 10906
rect 1996 10854 2026 10906
rect 2026 10854 2052 10906
rect 1756 10852 1812 10854
rect 1836 10852 1892 10854
rect 1916 10852 1972 10854
rect 1996 10852 2052 10854
rect 4756 10906 4812 10908
rect 4836 10906 4892 10908
rect 4916 10906 4972 10908
rect 4996 10906 5052 10908
rect 4756 10854 4782 10906
rect 4782 10854 4812 10906
rect 4836 10854 4846 10906
rect 4846 10854 4892 10906
rect 4916 10854 4962 10906
rect 4962 10854 4972 10906
rect 4996 10854 5026 10906
rect 5026 10854 5052 10906
rect 4756 10852 4812 10854
rect 4836 10852 4892 10854
rect 4916 10852 4972 10854
rect 4996 10852 5052 10854
rect 7756 10906 7812 10908
rect 7836 10906 7892 10908
rect 7916 10906 7972 10908
rect 7996 10906 8052 10908
rect 7756 10854 7782 10906
rect 7782 10854 7812 10906
rect 7836 10854 7846 10906
rect 7846 10854 7892 10906
rect 7916 10854 7962 10906
rect 7962 10854 7972 10906
rect 7996 10854 8026 10906
rect 8026 10854 8052 10906
rect 7756 10852 7812 10854
rect 7836 10852 7892 10854
rect 7916 10852 7972 10854
rect 7996 10852 8052 10854
rect 3256 10362 3312 10364
rect 3336 10362 3392 10364
rect 3416 10362 3472 10364
rect 3496 10362 3552 10364
rect 3256 10310 3282 10362
rect 3282 10310 3312 10362
rect 3336 10310 3346 10362
rect 3346 10310 3392 10362
rect 3416 10310 3462 10362
rect 3462 10310 3472 10362
rect 3496 10310 3526 10362
rect 3526 10310 3552 10362
rect 3256 10308 3312 10310
rect 3336 10308 3392 10310
rect 3416 10308 3472 10310
rect 3496 10308 3552 10310
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6416 10362 6472 10364
rect 6496 10362 6552 10364
rect 6256 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6416 10310 6462 10362
rect 6462 10310 6472 10362
rect 6496 10310 6526 10362
rect 6526 10310 6552 10362
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6416 10308 6472 10310
rect 6496 10308 6552 10310
rect 1756 9818 1812 9820
rect 1836 9818 1892 9820
rect 1916 9818 1972 9820
rect 1996 9818 2052 9820
rect 1756 9766 1782 9818
rect 1782 9766 1812 9818
rect 1836 9766 1846 9818
rect 1846 9766 1892 9818
rect 1916 9766 1962 9818
rect 1962 9766 1972 9818
rect 1996 9766 2026 9818
rect 2026 9766 2052 9818
rect 1756 9764 1812 9766
rect 1836 9764 1892 9766
rect 1916 9764 1972 9766
rect 1996 9764 2052 9766
rect 4756 9818 4812 9820
rect 4836 9818 4892 9820
rect 4916 9818 4972 9820
rect 4996 9818 5052 9820
rect 4756 9766 4782 9818
rect 4782 9766 4812 9818
rect 4836 9766 4846 9818
rect 4846 9766 4892 9818
rect 4916 9766 4962 9818
rect 4962 9766 4972 9818
rect 4996 9766 5026 9818
rect 5026 9766 5052 9818
rect 4756 9764 4812 9766
rect 4836 9764 4892 9766
rect 4916 9764 4972 9766
rect 4996 9764 5052 9766
rect 7756 9818 7812 9820
rect 7836 9818 7892 9820
rect 7916 9818 7972 9820
rect 7996 9818 8052 9820
rect 7756 9766 7782 9818
rect 7782 9766 7812 9818
rect 7836 9766 7846 9818
rect 7846 9766 7892 9818
rect 7916 9766 7962 9818
rect 7962 9766 7972 9818
rect 7996 9766 8026 9818
rect 8026 9766 8052 9818
rect 7756 9764 7812 9766
rect 7836 9764 7892 9766
rect 7916 9764 7972 9766
rect 7996 9764 8052 9766
rect 3256 9274 3312 9276
rect 3336 9274 3392 9276
rect 3416 9274 3472 9276
rect 3496 9274 3552 9276
rect 3256 9222 3282 9274
rect 3282 9222 3312 9274
rect 3336 9222 3346 9274
rect 3346 9222 3392 9274
rect 3416 9222 3462 9274
rect 3462 9222 3472 9274
rect 3496 9222 3526 9274
rect 3526 9222 3552 9274
rect 3256 9220 3312 9222
rect 3336 9220 3392 9222
rect 3416 9220 3472 9222
rect 3496 9220 3552 9222
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6416 9274 6472 9276
rect 6496 9274 6552 9276
rect 6256 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6416 9222 6462 9274
rect 6462 9222 6472 9274
rect 6496 9222 6526 9274
rect 6526 9222 6552 9274
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6416 9220 6472 9222
rect 6496 9220 6552 9222
rect 1756 8730 1812 8732
rect 1836 8730 1892 8732
rect 1916 8730 1972 8732
rect 1996 8730 2052 8732
rect 1756 8678 1782 8730
rect 1782 8678 1812 8730
rect 1836 8678 1846 8730
rect 1846 8678 1892 8730
rect 1916 8678 1962 8730
rect 1962 8678 1972 8730
rect 1996 8678 2026 8730
rect 2026 8678 2052 8730
rect 1756 8676 1812 8678
rect 1836 8676 1892 8678
rect 1916 8676 1972 8678
rect 1996 8676 2052 8678
rect 4756 8730 4812 8732
rect 4836 8730 4892 8732
rect 4916 8730 4972 8732
rect 4996 8730 5052 8732
rect 4756 8678 4782 8730
rect 4782 8678 4812 8730
rect 4836 8678 4846 8730
rect 4846 8678 4892 8730
rect 4916 8678 4962 8730
rect 4962 8678 4972 8730
rect 4996 8678 5026 8730
rect 5026 8678 5052 8730
rect 4756 8676 4812 8678
rect 4836 8676 4892 8678
rect 4916 8676 4972 8678
rect 4996 8676 5052 8678
rect 3256 8186 3312 8188
rect 3336 8186 3392 8188
rect 3416 8186 3472 8188
rect 3496 8186 3552 8188
rect 3256 8134 3282 8186
rect 3282 8134 3312 8186
rect 3336 8134 3346 8186
rect 3346 8134 3392 8186
rect 3416 8134 3462 8186
rect 3462 8134 3472 8186
rect 3496 8134 3526 8186
rect 3526 8134 3552 8186
rect 3256 8132 3312 8134
rect 3336 8132 3392 8134
rect 3416 8132 3472 8134
rect 3496 8132 3552 8134
rect 1756 7642 1812 7644
rect 1836 7642 1892 7644
rect 1916 7642 1972 7644
rect 1996 7642 2052 7644
rect 1756 7590 1782 7642
rect 1782 7590 1812 7642
rect 1836 7590 1846 7642
rect 1846 7590 1892 7642
rect 1916 7590 1962 7642
rect 1962 7590 1972 7642
rect 1996 7590 2026 7642
rect 2026 7590 2052 7642
rect 1756 7588 1812 7590
rect 1836 7588 1892 7590
rect 1916 7588 1972 7590
rect 1996 7588 2052 7590
rect 4756 7642 4812 7644
rect 4836 7642 4892 7644
rect 4916 7642 4972 7644
rect 4996 7642 5052 7644
rect 4756 7590 4782 7642
rect 4782 7590 4812 7642
rect 4836 7590 4846 7642
rect 4846 7590 4892 7642
rect 4916 7590 4962 7642
rect 4962 7590 4972 7642
rect 4996 7590 5026 7642
rect 5026 7590 5052 7642
rect 4756 7588 4812 7590
rect 4836 7588 4892 7590
rect 4916 7588 4972 7590
rect 4996 7588 5052 7590
rect 3256 7098 3312 7100
rect 3336 7098 3392 7100
rect 3416 7098 3472 7100
rect 3496 7098 3552 7100
rect 3256 7046 3282 7098
rect 3282 7046 3312 7098
rect 3336 7046 3346 7098
rect 3346 7046 3392 7098
rect 3416 7046 3462 7098
rect 3462 7046 3472 7098
rect 3496 7046 3526 7098
rect 3526 7046 3552 7098
rect 3256 7044 3312 7046
rect 3336 7044 3392 7046
rect 3416 7044 3472 7046
rect 3496 7044 3552 7046
rect 1756 6554 1812 6556
rect 1836 6554 1892 6556
rect 1916 6554 1972 6556
rect 1996 6554 2052 6556
rect 1756 6502 1782 6554
rect 1782 6502 1812 6554
rect 1836 6502 1846 6554
rect 1846 6502 1892 6554
rect 1916 6502 1962 6554
rect 1962 6502 1972 6554
rect 1996 6502 2026 6554
rect 2026 6502 2052 6554
rect 1756 6500 1812 6502
rect 1836 6500 1892 6502
rect 1916 6500 1972 6502
rect 1996 6500 2052 6502
rect 4756 6554 4812 6556
rect 4836 6554 4892 6556
rect 4916 6554 4972 6556
rect 4996 6554 5052 6556
rect 4756 6502 4782 6554
rect 4782 6502 4812 6554
rect 4836 6502 4846 6554
rect 4846 6502 4892 6554
rect 4916 6502 4962 6554
rect 4962 6502 4972 6554
rect 4996 6502 5026 6554
rect 5026 6502 5052 6554
rect 4756 6500 4812 6502
rect 4836 6500 4892 6502
rect 4916 6500 4972 6502
rect 4996 6500 5052 6502
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6416 8186 6472 8188
rect 6496 8186 6552 8188
rect 6256 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6416 8134 6462 8186
rect 6462 8134 6472 8186
rect 6496 8134 6526 8186
rect 6526 8134 6552 8186
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6416 8132 6472 8134
rect 6496 8132 6552 8134
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6416 7098 6472 7100
rect 6496 7098 6552 7100
rect 6256 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6416 7046 6462 7098
rect 6462 7046 6472 7098
rect 6496 7046 6526 7098
rect 6526 7046 6552 7098
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6416 7044 6472 7046
rect 6496 7044 6552 7046
rect 3256 6010 3312 6012
rect 3336 6010 3392 6012
rect 3416 6010 3472 6012
rect 3496 6010 3552 6012
rect 3256 5958 3282 6010
rect 3282 5958 3312 6010
rect 3336 5958 3346 6010
rect 3346 5958 3392 6010
rect 3416 5958 3462 6010
rect 3462 5958 3472 6010
rect 3496 5958 3526 6010
rect 3526 5958 3552 6010
rect 3256 5956 3312 5958
rect 3336 5956 3392 5958
rect 3416 5956 3472 5958
rect 3496 5956 3552 5958
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6416 6010 6472 6012
rect 6496 6010 6552 6012
rect 6256 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6416 5958 6462 6010
rect 6462 5958 6472 6010
rect 6496 5958 6526 6010
rect 6526 5958 6552 6010
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6416 5956 6472 5958
rect 6496 5956 6552 5958
rect 7756 8730 7812 8732
rect 7836 8730 7892 8732
rect 7916 8730 7972 8732
rect 7996 8730 8052 8732
rect 7756 8678 7782 8730
rect 7782 8678 7812 8730
rect 7836 8678 7846 8730
rect 7846 8678 7892 8730
rect 7916 8678 7962 8730
rect 7962 8678 7972 8730
rect 7996 8678 8026 8730
rect 8026 8678 8052 8730
rect 7756 8676 7812 8678
rect 7836 8676 7892 8678
rect 7916 8676 7972 8678
rect 7996 8676 8052 8678
rect 7756 7642 7812 7644
rect 7836 7642 7892 7644
rect 7916 7642 7972 7644
rect 7996 7642 8052 7644
rect 7756 7590 7782 7642
rect 7782 7590 7812 7642
rect 7836 7590 7846 7642
rect 7846 7590 7892 7642
rect 7916 7590 7962 7642
rect 7962 7590 7972 7642
rect 7996 7590 8026 7642
rect 8026 7590 8052 7642
rect 7756 7588 7812 7590
rect 7836 7588 7892 7590
rect 7916 7588 7972 7590
rect 7996 7588 8052 7590
rect 1756 5466 1812 5468
rect 1836 5466 1892 5468
rect 1916 5466 1972 5468
rect 1996 5466 2052 5468
rect 1756 5414 1782 5466
rect 1782 5414 1812 5466
rect 1836 5414 1846 5466
rect 1846 5414 1892 5466
rect 1916 5414 1962 5466
rect 1962 5414 1972 5466
rect 1996 5414 2026 5466
rect 2026 5414 2052 5466
rect 1756 5412 1812 5414
rect 1836 5412 1892 5414
rect 1916 5412 1972 5414
rect 1996 5412 2052 5414
rect 4756 5466 4812 5468
rect 4836 5466 4892 5468
rect 4916 5466 4972 5468
rect 4996 5466 5052 5468
rect 4756 5414 4782 5466
rect 4782 5414 4812 5466
rect 4836 5414 4846 5466
rect 4846 5414 4892 5466
rect 4916 5414 4962 5466
rect 4962 5414 4972 5466
rect 4996 5414 5026 5466
rect 5026 5414 5052 5466
rect 4756 5412 4812 5414
rect 4836 5412 4892 5414
rect 4916 5412 4972 5414
rect 4996 5412 5052 5414
rect 9256 13626 9312 13628
rect 9336 13626 9392 13628
rect 9416 13626 9472 13628
rect 9496 13626 9552 13628
rect 9256 13574 9282 13626
rect 9282 13574 9312 13626
rect 9336 13574 9346 13626
rect 9346 13574 9392 13626
rect 9416 13574 9462 13626
rect 9462 13574 9472 13626
rect 9496 13574 9526 13626
rect 9526 13574 9552 13626
rect 9256 13572 9312 13574
rect 9336 13572 9392 13574
rect 9416 13572 9472 13574
rect 9496 13572 9552 13574
rect 10756 13082 10812 13084
rect 10836 13082 10892 13084
rect 10916 13082 10972 13084
rect 10996 13082 11052 13084
rect 10756 13030 10782 13082
rect 10782 13030 10812 13082
rect 10836 13030 10846 13082
rect 10846 13030 10892 13082
rect 10916 13030 10962 13082
rect 10962 13030 10972 13082
rect 10996 13030 11026 13082
rect 11026 13030 11052 13082
rect 10756 13028 10812 13030
rect 10836 13028 10892 13030
rect 10916 13028 10972 13030
rect 10996 13028 11052 13030
rect 9256 12538 9312 12540
rect 9336 12538 9392 12540
rect 9416 12538 9472 12540
rect 9496 12538 9552 12540
rect 9256 12486 9282 12538
rect 9282 12486 9312 12538
rect 9336 12486 9346 12538
rect 9346 12486 9392 12538
rect 9416 12486 9462 12538
rect 9462 12486 9472 12538
rect 9496 12486 9526 12538
rect 9526 12486 9552 12538
rect 9256 12484 9312 12486
rect 9336 12484 9392 12486
rect 9416 12484 9472 12486
rect 9496 12484 9552 12486
rect 12256 13626 12312 13628
rect 12336 13626 12392 13628
rect 12416 13626 12472 13628
rect 12496 13626 12552 13628
rect 12256 13574 12282 13626
rect 12282 13574 12312 13626
rect 12336 13574 12346 13626
rect 12346 13574 12392 13626
rect 12416 13574 12462 13626
rect 12462 13574 12472 13626
rect 12496 13574 12526 13626
rect 12526 13574 12552 13626
rect 12256 13572 12312 13574
rect 12336 13572 12392 13574
rect 12416 13572 12472 13574
rect 12496 13572 12552 13574
rect 13756 15258 13812 15260
rect 13836 15258 13892 15260
rect 13916 15258 13972 15260
rect 13996 15258 14052 15260
rect 13756 15206 13782 15258
rect 13782 15206 13812 15258
rect 13836 15206 13846 15258
rect 13846 15206 13892 15258
rect 13916 15206 13962 15258
rect 13962 15206 13972 15258
rect 13996 15206 14026 15258
rect 14026 15206 14052 15258
rect 13756 15204 13812 15206
rect 13836 15204 13892 15206
rect 13916 15204 13972 15206
rect 13996 15204 14052 15206
rect 13756 14170 13812 14172
rect 13836 14170 13892 14172
rect 13916 14170 13972 14172
rect 13996 14170 14052 14172
rect 13756 14118 13782 14170
rect 13782 14118 13812 14170
rect 13836 14118 13846 14170
rect 13846 14118 13892 14170
rect 13916 14118 13962 14170
rect 13962 14118 13972 14170
rect 13996 14118 14026 14170
rect 14026 14118 14052 14170
rect 13756 14116 13812 14118
rect 13836 14116 13892 14118
rect 13916 14116 13972 14118
rect 13996 14116 14052 14118
rect 15256 15802 15312 15804
rect 15336 15802 15392 15804
rect 15416 15802 15472 15804
rect 15496 15802 15552 15804
rect 15256 15750 15282 15802
rect 15282 15750 15312 15802
rect 15336 15750 15346 15802
rect 15346 15750 15392 15802
rect 15416 15750 15462 15802
rect 15462 15750 15472 15802
rect 15496 15750 15526 15802
rect 15526 15750 15552 15802
rect 15256 15748 15312 15750
rect 15336 15748 15392 15750
rect 15416 15748 15472 15750
rect 15496 15748 15552 15750
rect 16756 16346 16812 16348
rect 16836 16346 16892 16348
rect 16916 16346 16972 16348
rect 16996 16346 17052 16348
rect 16756 16294 16782 16346
rect 16782 16294 16812 16346
rect 16836 16294 16846 16346
rect 16846 16294 16892 16346
rect 16916 16294 16962 16346
rect 16962 16294 16972 16346
rect 16996 16294 17026 16346
rect 17026 16294 17052 16346
rect 16756 16292 16812 16294
rect 16836 16292 16892 16294
rect 16916 16292 16972 16294
rect 16996 16292 17052 16294
rect 19756 16346 19812 16348
rect 19836 16346 19892 16348
rect 19916 16346 19972 16348
rect 19996 16346 20052 16348
rect 19756 16294 19782 16346
rect 19782 16294 19812 16346
rect 19836 16294 19846 16346
rect 19846 16294 19892 16346
rect 19916 16294 19962 16346
rect 19962 16294 19972 16346
rect 19996 16294 20026 16346
rect 20026 16294 20052 16346
rect 19756 16292 19812 16294
rect 19836 16292 19892 16294
rect 19916 16292 19972 16294
rect 19996 16292 20052 16294
rect 22756 16346 22812 16348
rect 22836 16346 22892 16348
rect 22916 16346 22972 16348
rect 22996 16346 23052 16348
rect 22756 16294 22782 16346
rect 22782 16294 22812 16346
rect 22836 16294 22846 16346
rect 22846 16294 22892 16346
rect 22916 16294 22962 16346
rect 22962 16294 22972 16346
rect 22996 16294 23026 16346
rect 23026 16294 23052 16346
rect 22756 16292 22812 16294
rect 22836 16292 22892 16294
rect 22916 16292 22972 16294
rect 22996 16292 23052 16294
rect 15256 14714 15312 14716
rect 15336 14714 15392 14716
rect 15416 14714 15472 14716
rect 15496 14714 15552 14716
rect 15256 14662 15282 14714
rect 15282 14662 15312 14714
rect 15336 14662 15346 14714
rect 15346 14662 15392 14714
rect 15416 14662 15462 14714
rect 15462 14662 15472 14714
rect 15496 14662 15526 14714
rect 15526 14662 15552 14714
rect 15256 14660 15312 14662
rect 15336 14660 15392 14662
rect 15416 14660 15472 14662
rect 15496 14660 15552 14662
rect 14278 14456 14334 14512
rect 14094 13912 14150 13968
rect 12256 12538 12312 12540
rect 12336 12538 12392 12540
rect 12416 12538 12472 12540
rect 12496 12538 12552 12540
rect 12256 12486 12282 12538
rect 12282 12486 12312 12538
rect 12336 12486 12346 12538
rect 12346 12486 12392 12538
rect 12416 12486 12462 12538
rect 12462 12486 12472 12538
rect 12496 12486 12526 12538
rect 12526 12486 12552 12538
rect 12256 12484 12312 12486
rect 12336 12484 12392 12486
rect 12416 12484 12472 12486
rect 12496 12484 12552 12486
rect 9256 11450 9312 11452
rect 9336 11450 9392 11452
rect 9416 11450 9472 11452
rect 9496 11450 9552 11452
rect 9256 11398 9282 11450
rect 9282 11398 9312 11450
rect 9336 11398 9346 11450
rect 9346 11398 9392 11450
rect 9416 11398 9462 11450
rect 9462 11398 9472 11450
rect 9496 11398 9526 11450
rect 9526 11398 9552 11450
rect 9256 11396 9312 11398
rect 9336 11396 9392 11398
rect 9416 11396 9472 11398
rect 9496 11396 9552 11398
rect 9256 10362 9312 10364
rect 9336 10362 9392 10364
rect 9416 10362 9472 10364
rect 9496 10362 9552 10364
rect 9256 10310 9282 10362
rect 9282 10310 9312 10362
rect 9336 10310 9346 10362
rect 9346 10310 9392 10362
rect 9416 10310 9462 10362
rect 9462 10310 9472 10362
rect 9496 10310 9526 10362
rect 9526 10310 9552 10362
rect 9256 10308 9312 10310
rect 9336 10308 9392 10310
rect 9416 10308 9472 10310
rect 9496 10308 9552 10310
rect 10756 11994 10812 11996
rect 10836 11994 10892 11996
rect 10916 11994 10972 11996
rect 10996 11994 11052 11996
rect 10756 11942 10782 11994
rect 10782 11942 10812 11994
rect 10836 11942 10846 11994
rect 10846 11942 10892 11994
rect 10916 11942 10962 11994
rect 10962 11942 10972 11994
rect 10996 11942 11026 11994
rect 11026 11942 11052 11994
rect 10756 11940 10812 11942
rect 10836 11940 10892 11942
rect 10916 11940 10972 11942
rect 10996 11940 11052 11942
rect 9256 9274 9312 9276
rect 9336 9274 9392 9276
rect 9416 9274 9472 9276
rect 9496 9274 9552 9276
rect 9256 9222 9282 9274
rect 9282 9222 9312 9274
rect 9336 9222 9346 9274
rect 9346 9222 9392 9274
rect 9416 9222 9462 9274
rect 9462 9222 9472 9274
rect 9496 9222 9526 9274
rect 9526 9222 9552 9274
rect 9256 9220 9312 9222
rect 9336 9220 9392 9222
rect 9416 9220 9472 9222
rect 9496 9220 9552 9222
rect 10756 10906 10812 10908
rect 10836 10906 10892 10908
rect 10916 10906 10972 10908
rect 10996 10906 11052 10908
rect 10756 10854 10782 10906
rect 10782 10854 10812 10906
rect 10836 10854 10846 10906
rect 10846 10854 10892 10906
rect 10916 10854 10962 10906
rect 10962 10854 10972 10906
rect 10996 10854 11026 10906
rect 11026 10854 11052 10906
rect 10756 10852 10812 10854
rect 10836 10852 10892 10854
rect 10916 10852 10972 10854
rect 10996 10852 11052 10854
rect 10756 9818 10812 9820
rect 10836 9818 10892 9820
rect 10916 9818 10972 9820
rect 10996 9818 11052 9820
rect 10756 9766 10782 9818
rect 10782 9766 10812 9818
rect 10836 9766 10846 9818
rect 10846 9766 10892 9818
rect 10916 9766 10962 9818
rect 10962 9766 10972 9818
rect 10996 9766 11026 9818
rect 11026 9766 11052 9818
rect 10756 9764 10812 9766
rect 10836 9764 10892 9766
rect 10916 9764 10972 9766
rect 10996 9764 11052 9766
rect 12256 11450 12312 11452
rect 12336 11450 12392 11452
rect 12416 11450 12472 11452
rect 12496 11450 12552 11452
rect 12256 11398 12282 11450
rect 12282 11398 12312 11450
rect 12336 11398 12346 11450
rect 12346 11398 12392 11450
rect 12416 11398 12462 11450
rect 12462 11398 12472 11450
rect 12496 11398 12526 11450
rect 12526 11398 12552 11450
rect 12256 11396 12312 11398
rect 12336 11396 12392 11398
rect 12416 11396 12472 11398
rect 12496 11396 12552 11398
rect 9256 8186 9312 8188
rect 9336 8186 9392 8188
rect 9416 8186 9472 8188
rect 9496 8186 9552 8188
rect 9256 8134 9282 8186
rect 9282 8134 9312 8186
rect 9336 8134 9346 8186
rect 9346 8134 9392 8186
rect 9416 8134 9462 8186
rect 9462 8134 9472 8186
rect 9496 8134 9526 8186
rect 9526 8134 9552 8186
rect 9256 8132 9312 8134
rect 9336 8132 9392 8134
rect 9416 8132 9472 8134
rect 9496 8132 9552 8134
rect 7756 6554 7812 6556
rect 7836 6554 7892 6556
rect 7916 6554 7972 6556
rect 7996 6554 8052 6556
rect 7756 6502 7782 6554
rect 7782 6502 7812 6554
rect 7836 6502 7846 6554
rect 7846 6502 7892 6554
rect 7916 6502 7962 6554
rect 7962 6502 7972 6554
rect 7996 6502 8026 6554
rect 8026 6502 8052 6554
rect 7756 6500 7812 6502
rect 7836 6500 7892 6502
rect 7916 6500 7972 6502
rect 7996 6500 8052 6502
rect 9256 7098 9312 7100
rect 9336 7098 9392 7100
rect 9416 7098 9472 7100
rect 9496 7098 9552 7100
rect 9256 7046 9282 7098
rect 9282 7046 9312 7098
rect 9336 7046 9346 7098
rect 9346 7046 9392 7098
rect 9416 7046 9462 7098
rect 9462 7046 9472 7098
rect 9496 7046 9526 7098
rect 9526 7046 9552 7098
rect 9256 7044 9312 7046
rect 9336 7044 9392 7046
rect 9416 7044 9472 7046
rect 9496 7044 9552 7046
rect 10756 8730 10812 8732
rect 10836 8730 10892 8732
rect 10916 8730 10972 8732
rect 10996 8730 11052 8732
rect 10756 8678 10782 8730
rect 10782 8678 10812 8730
rect 10836 8678 10846 8730
rect 10846 8678 10892 8730
rect 10916 8678 10962 8730
rect 10962 8678 10972 8730
rect 10996 8678 11026 8730
rect 11026 8678 11052 8730
rect 10756 8676 10812 8678
rect 10836 8676 10892 8678
rect 10916 8676 10972 8678
rect 10996 8676 11052 8678
rect 10756 7642 10812 7644
rect 10836 7642 10892 7644
rect 10916 7642 10972 7644
rect 10996 7642 11052 7644
rect 10756 7590 10782 7642
rect 10782 7590 10812 7642
rect 10836 7590 10846 7642
rect 10846 7590 10892 7642
rect 10916 7590 10962 7642
rect 10962 7590 10972 7642
rect 10996 7590 11026 7642
rect 11026 7590 11052 7642
rect 10756 7588 10812 7590
rect 10836 7588 10892 7590
rect 10916 7588 10972 7590
rect 10996 7588 11052 7590
rect 7756 5466 7812 5468
rect 7836 5466 7892 5468
rect 7916 5466 7972 5468
rect 7996 5466 8052 5468
rect 7756 5414 7782 5466
rect 7782 5414 7812 5466
rect 7836 5414 7846 5466
rect 7846 5414 7892 5466
rect 7916 5414 7962 5466
rect 7962 5414 7972 5466
rect 7996 5414 8026 5466
rect 8026 5414 8052 5466
rect 7756 5412 7812 5414
rect 7836 5412 7892 5414
rect 7916 5412 7972 5414
rect 7996 5412 8052 5414
rect 3256 4922 3312 4924
rect 3336 4922 3392 4924
rect 3416 4922 3472 4924
rect 3496 4922 3552 4924
rect 3256 4870 3282 4922
rect 3282 4870 3312 4922
rect 3336 4870 3346 4922
rect 3346 4870 3392 4922
rect 3416 4870 3462 4922
rect 3462 4870 3472 4922
rect 3496 4870 3526 4922
rect 3526 4870 3552 4922
rect 3256 4868 3312 4870
rect 3336 4868 3392 4870
rect 3416 4868 3472 4870
rect 3496 4868 3552 4870
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6416 4922 6472 4924
rect 6496 4922 6552 4924
rect 6256 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6416 4870 6462 4922
rect 6462 4870 6472 4922
rect 6496 4870 6526 4922
rect 6526 4870 6552 4922
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6416 4868 6472 4870
rect 6496 4868 6552 4870
rect 9256 6010 9312 6012
rect 9336 6010 9392 6012
rect 9416 6010 9472 6012
rect 9496 6010 9552 6012
rect 9256 5958 9282 6010
rect 9282 5958 9312 6010
rect 9336 5958 9346 6010
rect 9346 5958 9392 6010
rect 9416 5958 9462 6010
rect 9462 5958 9472 6010
rect 9496 5958 9526 6010
rect 9526 5958 9552 6010
rect 9256 5956 9312 5958
rect 9336 5956 9392 5958
rect 9416 5956 9472 5958
rect 9496 5956 9552 5958
rect 1756 4378 1812 4380
rect 1836 4378 1892 4380
rect 1916 4378 1972 4380
rect 1996 4378 2052 4380
rect 1756 4326 1782 4378
rect 1782 4326 1812 4378
rect 1836 4326 1846 4378
rect 1846 4326 1892 4378
rect 1916 4326 1962 4378
rect 1962 4326 1972 4378
rect 1996 4326 2026 4378
rect 2026 4326 2052 4378
rect 1756 4324 1812 4326
rect 1836 4324 1892 4326
rect 1916 4324 1972 4326
rect 1996 4324 2052 4326
rect 4756 4378 4812 4380
rect 4836 4378 4892 4380
rect 4916 4378 4972 4380
rect 4996 4378 5052 4380
rect 4756 4326 4782 4378
rect 4782 4326 4812 4378
rect 4836 4326 4846 4378
rect 4846 4326 4892 4378
rect 4916 4326 4962 4378
rect 4962 4326 4972 4378
rect 4996 4326 5026 4378
rect 5026 4326 5052 4378
rect 4756 4324 4812 4326
rect 4836 4324 4892 4326
rect 4916 4324 4972 4326
rect 4996 4324 5052 4326
rect 7756 4378 7812 4380
rect 7836 4378 7892 4380
rect 7916 4378 7972 4380
rect 7996 4378 8052 4380
rect 7756 4326 7782 4378
rect 7782 4326 7812 4378
rect 7836 4326 7846 4378
rect 7846 4326 7892 4378
rect 7916 4326 7962 4378
rect 7962 4326 7972 4378
rect 7996 4326 8026 4378
rect 8026 4326 8052 4378
rect 7756 4324 7812 4326
rect 7836 4324 7892 4326
rect 7916 4324 7972 4326
rect 7996 4324 8052 4326
rect 10756 6554 10812 6556
rect 10836 6554 10892 6556
rect 10916 6554 10972 6556
rect 10996 6554 11052 6556
rect 10756 6502 10782 6554
rect 10782 6502 10812 6554
rect 10836 6502 10846 6554
rect 10846 6502 10892 6554
rect 10916 6502 10962 6554
rect 10962 6502 10972 6554
rect 10996 6502 11026 6554
rect 11026 6502 11052 6554
rect 10756 6500 10812 6502
rect 10836 6500 10892 6502
rect 10916 6500 10972 6502
rect 10996 6500 11052 6502
rect 10756 5466 10812 5468
rect 10836 5466 10892 5468
rect 10916 5466 10972 5468
rect 10996 5466 11052 5468
rect 10756 5414 10782 5466
rect 10782 5414 10812 5466
rect 10836 5414 10846 5466
rect 10846 5414 10892 5466
rect 10916 5414 10962 5466
rect 10962 5414 10972 5466
rect 10996 5414 11026 5466
rect 11026 5414 11052 5466
rect 10756 5412 10812 5414
rect 10836 5412 10892 5414
rect 10916 5412 10972 5414
rect 10996 5412 11052 5414
rect 9256 4922 9312 4924
rect 9336 4922 9392 4924
rect 9416 4922 9472 4924
rect 9496 4922 9552 4924
rect 9256 4870 9282 4922
rect 9282 4870 9312 4922
rect 9336 4870 9346 4922
rect 9346 4870 9392 4922
rect 9416 4870 9462 4922
rect 9462 4870 9472 4922
rect 9496 4870 9526 4922
rect 9526 4870 9552 4922
rect 9256 4868 9312 4870
rect 9336 4868 9392 4870
rect 9416 4868 9472 4870
rect 9496 4868 9552 4870
rect 8850 4120 8906 4176
rect 3256 3834 3312 3836
rect 3336 3834 3392 3836
rect 3416 3834 3472 3836
rect 3496 3834 3552 3836
rect 3256 3782 3282 3834
rect 3282 3782 3312 3834
rect 3336 3782 3346 3834
rect 3346 3782 3392 3834
rect 3416 3782 3462 3834
rect 3462 3782 3472 3834
rect 3496 3782 3526 3834
rect 3526 3782 3552 3834
rect 3256 3780 3312 3782
rect 3336 3780 3392 3782
rect 3416 3780 3472 3782
rect 3496 3780 3552 3782
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6416 3834 6472 3836
rect 6496 3834 6552 3836
rect 6256 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6416 3782 6462 3834
rect 6462 3782 6472 3834
rect 6496 3782 6526 3834
rect 6526 3782 6552 3834
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6416 3780 6472 3782
rect 6496 3780 6552 3782
rect 1756 3290 1812 3292
rect 1836 3290 1892 3292
rect 1916 3290 1972 3292
rect 1996 3290 2052 3292
rect 1756 3238 1782 3290
rect 1782 3238 1812 3290
rect 1836 3238 1846 3290
rect 1846 3238 1892 3290
rect 1916 3238 1962 3290
rect 1962 3238 1972 3290
rect 1996 3238 2026 3290
rect 2026 3238 2052 3290
rect 1756 3236 1812 3238
rect 1836 3236 1892 3238
rect 1916 3236 1972 3238
rect 1996 3236 2052 3238
rect 4756 3290 4812 3292
rect 4836 3290 4892 3292
rect 4916 3290 4972 3292
rect 4996 3290 5052 3292
rect 4756 3238 4782 3290
rect 4782 3238 4812 3290
rect 4836 3238 4846 3290
rect 4846 3238 4892 3290
rect 4916 3238 4962 3290
rect 4962 3238 4972 3290
rect 4996 3238 5026 3290
rect 5026 3238 5052 3290
rect 4756 3236 4812 3238
rect 4836 3236 4892 3238
rect 4916 3236 4972 3238
rect 4996 3236 5052 3238
rect 7756 3290 7812 3292
rect 7836 3290 7892 3292
rect 7916 3290 7972 3292
rect 7996 3290 8052 3292
rect 7756 3238 7782 3290
rect 7782 3238 7812 3290
rect 7836 3238 7846 3290
rect 7846 3238 7892 3290
rect 7916 3238 7962 3290
rect 7962 3238 7972 3290
rect 7996 3238 8026 3290
rect 8026 3238 8052 3290
rect 7756 3236 7812 3238
rect 7836 3236 7892 3238
rect 7916 3236 7972 3238
rect 7996 3236 8052 3238
rect 8758 3984 8814 4040
rect 3256 2746 3312 2748
rect 3336 2746 3392 2748
rect 3416 2746 3472 2748
rect 3496 2746 3552 2748
rect 3256 2694 3282 2746
rect 3282 2694 3312 2746
rect 3336 2694 3346 2746
rect 3346 2694 3392 2746
rect 3416 2694 3462 2746
rect 3462 2694 3472 2746
rect 3496 2694 3526 2746
rect 3526 2694 3552 2746
rect 3256 2692 3312 2694
rect 3336 2692 3392 2694
rect 3416 2692 3472 2694
rect 3496 2692 3552 2694
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6416 2746 6472 2748
rect 6496 2746 6552 2748
rect 6256 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6416 2694 6462 2746
rect 6462 2694 6472 2746
rect 6496 2694 6526 2746
rect 6526 2694 6552 2746
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 6416 2692 6472 2694
rect 6496 2692 6552 2694
rect 9256 3834 9312 3836
rect 9336 3834 9392 3836
rect 9416 3834 9472 3836
rect 9496 3834 9552 3836
rect 9256 3782 9282 3834
rect 9282 3782 9312 3834
rect 9336 3782 9346 3834
rect 9346 3782 9392 3834
rect 9416 3782 9462 3834
rect 9462 3782 9472 3834
rect 9496 3782 9526 3834
rect 9526 3782 9552 3834
rect 9256 3780 9312 3782
rect 9336 3780 9392 3782
rect 9416 3780 9472 3782
rect 9496 3780 9552 3782
rect 9954 3984 10010 4040
rect 1756 2202 1812 2204
rect 1836 2202 1892 2204
rect 1916 2202 1972 2204
rect 1996 2202 2052 2204
rect 1756 2150 1782 2202
rect 1782 2150 1812 2202
rect 1836 2150 1846 2202
rect 1846 2150 1892 2202
rect 1916 2150 1962 2202
rect 1962 2150 1972 2202
rect 1996 2150 2026 2202
rect 2026 2150 2052 2202
rect 1756 2148 1812 2150
rect 1836 2148 1892 2150
rect 1916 2148 1972 2150
rect 1996 2148 2052 2150
rect 4756 2202 4812 2204
rect 4836 2202 4892 2204
rect 4916 2202 4972 2204
rect 4996 2202 5052 2204
rect 4756 2150 4782 2202
rect 4782 2150 4812 2202
rect 4836 2150 4846 2202
rect 4846 2150 4892 2202
rect 4916 2150 4962 2202
rect 4962 2150 4972 2202
rect 4996 2150 5026 2202
rect 5026 2150 5052 2202
rect 4756 2148 4812 2150
rect 4836 2148 4892 2150
rect 4916 2148 4972 2150
rect 4996 2148 5052 2150
rect 7756 2202 7812 2204
rect 7836 2202 7892 2204
rect 7916 2202 7972 2204
rect 7996 2202 8052 2204
rect 7756 2150 7782 2202
rect 7782 2150 7812 2202
rect 7836 2150 7846 2202
rect 7846 2150 7892 2202
rect 7916 2150 7962 2202
rect 7962 2150 7972 2202
rect 7996 2150 8026 2202
rect 8026 2150 8052 2202
rect 7756 2148 7812 2150
rect 7836 2148 7892 2150
rect 7916 2148 7972 2150
rect 7996 2148 8052 2150
rect 9256 2746 9312 2748
rect 9336 2746 9392 2748
rect 9416 2746 9472 2748
rect 9496 2746 9552 2748
rect 9256 2694 9282 2746
rect 9282 2694 9312 2746
rect 9336 2694 9346 2746
rect 9346 2694 9392 2746
rect 9416 2694 9462 2746
rect 9462 2694 9472 2746
rect 9496 2694 9526 2746
rect 9526 2694 9552 2746
rect 9256 2692 9312 2694
rect 9336 2692 9392 2694
rect 9416 2692 9472 2694
rect 9496 2692 9552 2694
rect 10756 4378 10812 4380
rect 10836 4378 10892 4380
rect 10916 4378 10972 4380
rect 10996 4378 11052 4380
rect 10756 4326 10782 4378
rect 10782 4326 10812 4378
rect 10836 4326 10846 4378
rect 10846 4326 10892 4378
rect 10916 4326 10962 4378
rect 10962 4326 10972 4378
rect 10996 4326 11026 4378
rect 11026 4326 11052 4378
rect 10756 4324 10812 4326
rect 10836 4324 10892 4326
rect 10916 4324 10972 4326
rect 10996 4324 11052 4326
rect 10756 3290 10812 3292
rect 10836 3290 10892 3292
rect 10916 3290 10972 3292
rect 10996 3290 11052 3292
rect 10756 3238 10782 3290
rect 10782 3238 10812 3290
rect 10836 3238 10846 3290
rect 10846 3238 10892 3290
rect 10916 3238 10962 3290
rect 10962 3238 10972 3290
rect 10996 3238 11026 3290
rect 11026 3238 11052 3290
rect 10756 3236 10812 3238
rect 10836 3236 10892 3238
rect 10916 3236 10972 3238
rect 10996 3236 11052 3238
rect 15256 13626 15312 13628
rect 15336 13626 15392 13628
rect 15416 13626 15472 13628
rect 15496 13626 15552 13628
rect 15256 13574 15282 13626
rect 15282 13574 15312 13626
rect 15336 13574 15346 13626
rect 15346 13574 15392 13626
rect 15416 13574 15462 13626
rect 15462 13574 15472 13626
rect 15496 13574 15526 13626
rect 15526 13574 15552 13626
rect 15256 13572 15312 13574
rect 15336 13572 15392 13574
rect 15416 13572 15472 13574
rect 15496 13572 15552 13574
rect 16756 15258 16812 15260
rect 16836 15258 16892 15260
rect 16916 15258 16972 15260
rect 16996 15258 17052 15260
rect 16756 15206 16782 15258
rect 16782 15206 16812 15258
rect 16836 15206 16846 15258
rect 16846 15206 16892 15258
rect 16916 15206 16962 15258
rect 16962 15206 16972 15258
rect 16996 15206 17026 15258
rect 17026 15206 17052 15258
rect 16756 15204 16812 15206
rect 16836 15204 16892 15206
rect 16916 15204 16972 15206
rect 16996 15204 17052 15206
rect 18256 15802 18312 15804
rect 18336 15802 18392 15804
rect 18416 15802 18472 15804
rect 18496 15802 18552 15804
rect 18256 15750 18282 15802
rect 18282 15750 18312 15802
rect 18336 15750 18346 15802
rect 18346 15750 18392 15802
rect 18416 15750 18462 15802
rect 18462 15750 18472 15802
rect 18496 15750 18526 15802
rect 18526 15750 18552 15802
rect 18256 15748 18312 15750
rect 18336 15748 18392 15750
rect 18416 15748 18472 15750
rect 18496 15748 18552 15750
rect 13756 13082 13812 13084
rect 13836 13082 13892 13084
rect 13916 13082 13972 13084
rect 13996 13082 14052 13084
rect 13756 13030 13782 13082
rect 13782 13030 13812 13082
rect 13836 13030 13846 13082
rect 13846 13030 13892 13082
rect 13916 13030 13962 13082
rect 13962 13030 13972 13082
rect 13996 13030 14026 13082
rect 14026 13030 14052 13082
rect 13756 13028 13812 13030
rect 13836 13028 13892 13030
rect 13916 13028 13972 13030
rect 13996 13028 14052 13030
rect 13756 11994 13812 11996
rect 13836 11994 13892 11996
rect 13916 11994 13972 11996
rect 13996 11994 14052 11996
rect 13756 11942 13782 11994
rect 13782 11942 13812 11994
rect 13836 11942 13846 11994
rect 13846 11942 13892 11994
rect 13916 11942 13962 11994
rect 13962 11942 13972 11994
rect 13996 11942 14026 11994
rect 14026 11942 14052 11994
rect 13756 11940 13812 11942
rect 13836 11940 13892 11942
rect 13916 11940 13972 11942
rect 13996 11940 14052 11942
rect 13756 10906 13812 10908
rect 13836 10906 13892 10908
rect 13916 10906 13972 10908
rect 13996 10906 14052 10908
rect 13756 10854 13782 10906
rect 13782 10854 13812 10906
rect 13836 10854 13846 10906
rect 13846 10854 13892 10906
rect 13916 10854 13962 10906
rect 13962 10854 13972 10906
rect 13996 10854 14026 10906
rect 14026 10854 14052 10906
rect 13756 10852 13812 10854
rect 13836 10852 13892 10854
rect 13916 10852 13972 10854
rect 13996 10852 14052 10854
rect 12256 10362 12312 10364
rect 12336 10362 12392 10364
rect 12416 10362 12472 10364
rect 12496 10362 12552 10364
rect 12256 10310 12282 10362
rect 12282 10310 12312 10362
rect 12336 10310 12346 10362
rect 12346 10310 12392 10362
rect 12416 10310 12462 10362
rect 12462 10310 12472 10362
rect 12496 10310 12526 10362
rect 12526 10310 12552 10362
rect 12256 10308 12312 10310
rect 12336 10308 12392 10310
rect 12416 10308 12472 10310
rect 12496 10308 12552 10310
rect 12256 9274 12312 9276
rect 12336 9274 12392 9276
rect 12416 9274 12472 9276
rect 12496 9274 12552 9276
rect 12256 9222 12282 9274
rect 12282 9222 12312 9274
rect 12336 9222 12346 9274
rect 12346 9222 12392 9274
rect 12416 9222 12462 9274
rect 12462 9222 12472 9274
rect 12496 9222 12526 9274
rect 12526 9222 12552 9274
rect 12256 9220 12312 9222
rect 12336 9220 12392 9222
rect 12416 9220 12472 9222
rect 12496 9220 12552 9222
rect 13756 9818 13812 9820
rect 13836 9818 13892 9820
rect 13916 9818 13972 9820
rect 13996 9818 14052 9820
rect 13756 9766 13782 9818
rect 13782 9766 13812 9818
rect 13836 9766 13846 9818
rect 13846 9766 13892 9818
rect 13916 9766 13962 9818
rect 13962 9766 13972 9818
rect 13996 9766 14026 9818
rect 14026 9766 14052 9818
rect 13756 9764 13812 9766
rect 13836 9764 13892 9766
rect 13916 9764 13972 9766
rect 13996 9764 14052 9766
rect 13756 8730 13812 8732
rect 13836 8730 13892 8732
rect 13916 8730 13972 8732
rect 13996 8730 14052 8732
rect 13756 8678 13782 8730
rect 13782 8678 13812 8730
rect 13836 8678 13846 8730
rect 13846 8678 13892 8730
rect 13916 8678 13962 8730
rect 13962 8678 13972 8730
rect 13996 8678 14026 8730
rect 14026 8678 14052 8730
rect 13756 8676 13812 8678
rect 13836 8676 13892 8678
rect 13916 8676 13972 8678
rect 13996 8676 14052 8678
rect 12256 8186 12312 8188
rect 12336 8186 12392 8188
rect 12416 8186 12472 8188
rect 12496 8186 12552 8188
rect 12256 8134 12282 8186
rect 12282 8134 12312 8186
rect 12336 8134 12346 8186
rect 12346 8134 12392 8186
rect 12416 8134 12462 8186
rect 12462 8134 12472 8186
rect 12496 8134 12526 8186
rect 12526 8134 12552 8186
rect 12256 8132 12312 8134
rect 12336 8132 12392 8134
rect 12416 8132 12472 8134
rect 12496 8132 12552 8134
rect 13756 7642 13812 7644
rect 13836 7642 13892 7644
rect 13916 7642 13972 7644
rect 13996 7642 14052 7644
rect 13756 7590 13782 7642
rect 13782 7590 13812 7642
rect 13836 7590 13846 7642
rect 13846 7590 13892 7642
rect 13916 7590 13962 7642
rect 13962 7590 13972 7642
rect 13996 7590 14026 7642
rect 14026 7590 14052 7642
rect 13756 7588 13812 7590
rect 13836 7588 13892 7590
rect 13916 7588 13972 7590
rect 13996 7588 14052 7590
rect 11794 4120 11850 4176
rect 12256 7098 12312 7100
rect 12336 7098 12392 7100
rect 12416 7098 12472 7100
rect 12496 7098 12552 7100
rect 12256 7046 12282 7098
rect 12282 7046 12312 7098
rect 12336 7046 12346 7098
rect 12346 7046 12392 7098
rect 12416 7046 12462 7098
rect 12462 7046 12472 7098
rect 12496 7046 12526 7098
rect 12526 7046 12552 7098
rect 12256 7044 12312 7046
rect 12336 7044 12392 7046
rect 12416 7044 12472 7046
rect 12496 7044 12552 7046
rect 12256 6010 12312 6012
rect 12336 6010 12392 6012
rect 12416 6010 12472 6012
rect 12496 6010 12552 6012
rect 12256 5958 12282 6010
rect 12282 5958 12312 6010
rect 12336 5958 12346 6010
rect 12346 5958 12392 6010
rect 12416 5958 12462 6010
rect 12462 5958 12472 6010
rect 12496 5958 12526 6010
rect 12526 5958 12552 6010
rect 12256 5956 12312 5958
rect 12336 5956 12392 5958
rect 12416 5956 12472 5958
rect 12496 5956 12552 5958
rect 13756 6554 13812 6556
rect 13836 6554 13892 6556
rect 13916 6554 13972 6556
rect 13996 6554 14052 6556
rect 13756 6502 13782 6554
rect 13782 6502 13812 6554
rect 13836 6502 13846 6554
rect 13846 6502 13892 6554
rect 13916 6502 13962 6554
rect 13962 6502 13972 6554
rect 13996 6502 14026 6554
rect 14026 6502 14052 6554
rect 13756 6500 13812 6502
rect 13836 6500 13892 6502
rect 13916 6500 13972 6502
rect 13996 6500 14052 6502
rect 12070 4120 12126 4176
rect 12256 4922 12312 4924
rect 12336 4922 12392 4924
rect 12416 4922 12472 4924
rect 12496 4922 12552 4924
rect 12256 4870 12282 4922
rect 12282 4870 12312 4922
rect 12336 4870 12346 4922
rect 12346 4870 12392 4922
rect 12416 4870 12462 4922
rect 12462 4870 12472 4922
rect 12496 4870 12526 4922
rect 12526 4870 12552 4922
rect 12256 4868 12312 4870
rect 12336 4868 12392 4870
rect 12416 4868 12472 4870
rect 12496 4868 12552 4870
rect 12256 3834 12312 3836
rect 12336 3834 12392 3836
rect 12416 3834 12472 3836
rect 12496 3834 12552 3836
rect 12256 3782 12282 3834
rect 12282 3782 12312 3834
rect 12336 3782 12346 3834
rect 12346 3782 12392 3834
rect 12416 3782 12462 3834
rect 12462 3782 12472 3834
rect 12496 3782 12526 3834
rect 12526 3782 12552 3834
rect 12256 3780 12312 3782
rect 12336 3780 12392 3782
rect 12416 3780 12472 3782
rect 12496 3780 12552 3782
rect 13756 5466 13812 5468
rect 13836 5466 13892 5468
rect 13916 5466 13972 5468
rect 13996 5466 14052 5468
rect 13756 5414 13782 5466
rect 13782 5414 13812 5466
rect 13836 5414 13846 5466
rect 13846 5414 13892 5466
rect 13916 5414 13962 5466
rect 13962 5414 13972 5466
rect 13996 5414 14026 5466
rect 14026 5414 14052 5466
rect 13756 5412 13812 5414
rect 13836 5412 13892 5414
rect 13916 5412 13972 5414
rect 13996 5412 14052 5414
rect 13756 4378 13812 4380
rect 13836 4378 13892 4380
rect 13916 4378 13972 4380
rect 13996 4378 14052 4380
rect 13756 4326 13782 4378
rect 13782 4326 13812 4378
rect 13836 4326 13846 4378
rect 13846 4326 13892 4378
rect 13916 4326 13962 4378
rect 13962 4326 13972 4378
rect 13996 4326 14026 4378
rect 14026 4326 14052 4378
rect 13756 4324 13812 4326
rect 13836 4324 13892 4326
rect 13916 4324 13972 4326
rect 13996 4324 14052 4326
rect 15256 12538 15312 12540
rect 15336 12538 15392 12540
rect 15416 12538 15472 12540
rect 15496 12538 15552 12540
rect 15256 12486 15282 12538
rect 15282 12486 15312 12538
rect 15336 12486 15346 12538
rect 15346 12486 15392 12538
rect 15416 12486 15462 12538
rect 15462 12486 15472 12538
rect 15496 12486 15526 12538
rect 15526 12486 15552 12538
rect 15256 12484 15312 12486
rect 15336 12484 15392 12486
rect 15416 12484 15472 12486
rect 15496 12484 15552 12486
rect 15256 11450 15312 11452
rect 15336 11450 15392 11452
rect 15416 11450 15472 11452
rect 15496 11450 15552 11452
rect 15256 11398 15282 11450
rect 15282 11398 15312 11450
rect 15336 11398 15346 11450
rect 15346 11398 15392 11450
rect 15416 11398 15462 11450
rect 15462 11398 15472 11450
rect 15496 11398 15526 11450
rect 15526 11398 15552 11450
rect 15256 11396 15312 11398
rect 15336 11396 15392 11398
rect 15416 11396 15472 11398
rect 15496 11396 15552 11398
rect 15256 10362 15312 10364
rect 15336 10362 15392 10364
rect 15416 10362 15472 10364
rect 15496 10362 15552 10364
rect 15256 10310 15282 10362
rect 15282 10310 15312 10362
rect 15336 10310 15346 10362
rect 15346 10310 15392 10362
rect 15416 10310 15462 10362
rect 15462 10310 15472 10362
rect 15496 10310 15526 10362
rect 15526 10310 15552 10362
rect 15256 10308 15312 10310
rect 15336 10308 15392 10310
rect 15416 10308 15472 10310
rect 15496 10308 15552 10310
rect 15256 9274 15312 9276
rect 15336 9274 15392 9276
rect 15416 9274 15472 9276
rect 15496 9274 15552 9276
rect 15256 9222 15282 9274
rect 15282 9222 15312 9274
rect 15336 9222 15346 9274
rect 15346 9222 15392 9274
rect 15416 9222 15462 9274
rect 15462 9222 15472 9274
rect 15496 9222 15526 9274
rect 15526 9222 15552 9274
rect 15256 9220 15312 9222
rect 15336 9220 15392 9222
rect 15416 9220 15472 9222
rect 15496 9220 15552 9222
rect 15256 8186 15312 8188
rect 15336 8186 15392 8188
rect 15416 8186 15472 8188
rect 15496 8186 15552 8188
rect 15256 8134 15282 8186
rect 15282 8134 15312 8186
rect 15336 8134 15346 8186
rect 15346 8134 15392 8186
rect 15416 8134 15462 8186
rect 15462 8134 15472 8186
rect 15496 8134 15526 8186
rect 15526 8134 15552 8186
rect 15256 8132 15312 8134
rect 15336 8132 15392 8134
rect 15416 8132 15472 8134
rect 15496 8132 15552 8134
rect 15256 7098 15312 7100
rect 15336 7098 15392 7100
rect 15416 7098 15472 7100
rect 15496 7098 15552 7100
rect 15256 7046 15282 7098
rect 15282 7046 15312 7098
rect 15336 7046 15346 7098
rect 15346 7046 15392 7098
rect 15416 7046 15462 7098
rect 15462 7046 15472 7098
rect 15496 7046 15526 7098
rect 15526 7046 15552 7098
rect 15256 7044 15312 7046
rect 15336 7044 15392 7046
rect 15416 7044 15472 7046
rect 15496 7044 15552 7046
rect 12256 2746 12312 2748
rect 12336 2746 12392 2748
rect 12416 2746 12472 2748
rect 12496 2746 12552 2748
rect 12256 2694 12282 2746
rect 12282 2694 12312 2746
rect 12336 2694 12346 2746
rect 12346 2694 12392 2746
rect 12416 2694 12462 2746
rect 12462 2694 12472 2746
rect 12496 2694 12526 2746
rect 12526 2694 12552 2746
rect 12256 2692 12312 2694
rect 12336 2692 12392 2694
rect 12416 2692 12472 2694
rect 12496 2692 12552 2694
rect 13756 3290 13812 3292
rect 13836 3290 13892 3292
rect 13916 3290 13972 3292
rect 13996 3290 14052 3292
rect 13756 3238 13782 3290
rect 13782 3238 13812 3290
rect 13836 3238 13846 3290
rect 13846 3238 13892 3290
rect 13916 3238 13962 3290
rect 13962 3238 13972 3290
rect 13996 3238 14026 3290
rect 14026 3238 14052 3290
rect 13756 3236 13812 3238
rect 13836 3236 13892 3238
rect 13916 3236 13972 3238
rect 13996 3236 14052 3238
rect 15256 6010 15312 6012
rect 15336 6010 15392 6012
rect 15416 6010 15472 6012
rect 15496 6010 15552 6012
rect 15256 5958 15282 6010
rect 15282 5958 15312 6010
rect 15336 5958 15346 6010
rect 15346 5958 15392 6010
rect 15416 5958 15462 6010
rect 15462 5958 15472 6010
rect 15496 5958 15526 6010
rect 15526 5958 15552 6010
rect 15256 5956 15312 5958
rect 15336 5956 15392 5958
rect 15416 5956 15472 5958
rect 15496 5956 15552 5958
rect 16756 14170 16812 14172
rect 16836 14170 16892 14172
rect 16916 14170 16972 14172
rect 16996 14170 17052 14172
rect 16756 14118 16782 14170
rect 16782 14118 16812 14170
rect 16836 14118 16846 14170
rect 16846 14118 16892 14170
rect 16916 14118 16962 14170
rect 16962 14118 16972 14170
rect 16996 14118 17026 14170
rect 17026 14118 17052 14170
rect 16756 14116 16812 14118
rect 16836 14116 16892 14118
rect 16916 14116 16972 14118
rect 16996 14116 17052 14118
rect 16756 13082 16812 13084
rect 16836 13082 16892 13084
rect 16916 13082 16972 13084
rect 16996 13082 17052 13084
rect 16756 13030 16782 13082
rect 16782 13030 16812 13082
rect 16836 13030 16846 13082
rect 16846 13030 16892 13082
rect 16916 13030 16962 13082
rect 16962 13030 16972 13082
rect 16996 13030 17026 13082
rect 17026 13030 17052 13082
rect 16756 13028 16812 13030
rect 16836 13028 16892 13030
rect 16916 13028 16972 13030
rect 16996 13028 17052 13030
rect 16756 11994 16812 11996
rect 16836 11994 16892 11996
rect 16916 11994 16972 11996
rect 16996 11994 17052 11996
rect 16756 11942 16782 11994
rect 16782 11942 16812 11994
rect 16836 11942 16846 11994
rect 16846 11942 16892 11994
rect 16916 11942 16962 11994
rect 16962 11942 16972 11994
rect 16996 11942 17026 11994
rect 17026 11942 17052 11994
rect 16756 11940 16812 11942
rect 16836 11940 16892 11942
rect 16916 11940 16972 11942
rect 16996 11940 17052 11942
rect 18256 14714 18312 14716
rect 18336 14714 18392 14716
rect 18416 14714 18472 14716
rect 18496 14714 18552 14716
rect 18256 14662 18282 14714
rect 18282 14662 18312 14714
rect 18336 14662 18346 14714
rect 18346 14662 18392 14714
rect 18416 14662 18462 14714
rect 18462 14662 18472 14714
rect 18496 14662 18526 14714
rect 18526 14662 18552 14714
rect 18256 14660 18312 14662
rect 18336 14660 18392 14662
rect 18416 14660 18472 14662
rect 18496 14660 18552 14662
rect 16756 10906 16812 10908
rect 16836 10906 16892 10908
rect 16916 10906 16972 10908
rect 16996 10906 17052 10908
rect 16756 10854 16782 10906
rect 16782 10854 16812 10906
rect 16836 10854 16846 10906
rect 16846 10854 16892 10906
rect 16916 10854 16962 10906
rect 16962 10854 16972 10906
rect 16996 10854 17026 10906
rect 17026 10854 17052 10906
rect 16756 10852 16812 10854
rect 16836 10852 16892 10854
rect 16916 10852 16972 10854
rect 16996 10852 17052 10854
rect 15256 4922 15312 4924
rect 15336 4922 15392 4924
rect 15416 4922 15472 4924
rect 15496 4922 15552 4924
rect 15256 4870 15282 4922
rect 15282 4870 15312 4922
rect 15336 4870 15346 4922
rect 15346 4870 15392 4922
rect 15416 4870 15462 4922
rect 15462 4870 15472 4922
rect 15496 4870 15526 4922
rect 15526 4870 15552 4922
rect 15256 4868 15312 4870
rect 15336 4868 15392 4870
rect 15416 4868 15472 4870
rect 15496 4868 15552 4870
rect 15256 3834 15312 3836
rect 15336 3834 15392 3836
rect 15416 3834 15472 3836
rect 15496 3834 15552 3836
rect 15256 3782 15282 3834
rect 15282 3782 15312 3834
rect 15336 3782 15346 3834
rect 15346 3782 15392 3834
rect 15416 3782 15462 3834
rect 15462 3782 15472 3834
rect 15496 3782 15526 3834
rect 15526 3782 15552 3834
rect 15256 3780 15312 3782
rect 15336 3780 15392 3782
rect 15416 3780 15472 3782
rect 15496 3780 15552 3782
rect 16756 9818 16812 9820
rect 16836 9818 16892 9820
rect 16916 9818 16972 9820
rect 16996 9818 17052 9820
rect 16756 9766 16782 9818
rect 16782 9766 16812 9818
rect 16836 9766 16846 9818
rect 16846 9766 16892 9818
rect 16916 9766 16962 9818
rect 16962 9766 16972 9818
rect 16996 9766 17026 9818
rect 17026 9766 17052 9818
rect 16756 9764 16812 9766
rect 16836 9764 16892 9766
rect 16916 9764 16972 9766
rect 16996 9764 17052 9766
rect 18256 13626 18312 13628
rect 18336 13626 18392 13628
rect 18416 13626 18472 13628
rect 18496 13626 18552 13628
rect 18256 13574 18282 13626
rect 18282 13574 18312 13626
rect 18336 13574 18346 13626
rect 18346 13574 18392 13626
rect 18416 13574 18462 13626
rect 18462 13574 18472 13626
rect 18496 13574 18526 13626
rect 18526 13574 18552 13626
rect 18256 13572 18312 13574
rect 18336 13572 18392 13574
rect 18416 13572 18472 13574
rect 18496 13572 18552 13574
rect 18256 12538 18312 12540
rect 18336 12538 18392 12540
rect 18416 12538 18472 12540
rect 18496 12538 18552 12540
rect 18256 12486 18282 12538
rect 18282 12486 18312 12538
rect 18336 12486 18346 12538
rect 18346 12486 18392 12538
rect 18416 12486 18462 12538
rect 18462 12486 18472 12538
rect 18496 12486 18526 12538
rect 18526 12486 18552 12538
rect 18256 12484 18312 12486
rect 18336 12484 18392 12486
rect 18416 12484 18472 12486
rect 18496 12484 18552 12486
rect 21256 15802 21312 15804
rect 21336 15802 21392 15804
rect 21416 15802 21472 15804
rect 21496 15802 21552 15804
rect 21256 15750 21282 15802
rect 21282 15750 21312 15802
rect 21336 15750 21346 15802
rect 21346 15750 21392 15802
rect 21416 15750 21462 15802
rect 21462 15750 21472 15802
rect 21496 15750 21526 15802
rect 21526 15750 21552 15802
rect 21256 15748 21312 15750
rect 21336 15748 21392 15750
rect 21416 15748 21472 15750
rect 21496 15748 21552 15750
rect 19756 15258 19812 15260
rect 19836 15258 19892 15260
rect 19916 15258 19972 15260
rect 19996 15258 20052 15260
rect 19756 15206 19782 15258
rect 19782 15206 19812 15258
rect 19836 15206 19846 15258
rect 19846 15206 19892 15258
rect 19916 15206 19962 15258
rect 19962 15206 19972 15258
rect 19996 15206 20026 15258
rect 20026 15206 20052 15258
rect 19756 15204 19812 15206
rect 19836 15204 19892 15206
rect 19916 15204 19972 15206
rect 19996 15204 20052 15206
rect 19756 14170 19812 14172
rect 19836 14170 19892 14172
rect 19916 14170 19972 14172
rect 19996 14170 20052 14172
rect 19756 14118 19782 14170
rect 19782 14118 19812 14170
rect 19836 14118 19846 14170
rect 19846 14118 19892 14170
rect 19916 14118 19962 14170
rect 19962 14118 19972 14170
rect 19996 14118 20026 14170
rect 20026 14118 20052 14170
rect 19756 14116 19812 14118
rect 19836 14116 19892 14118
rect 19916 14116 19972 14118
rect 19996 14116 20052 14118
rect 19756 13082 19812 13084
rect 19836 13082 19892 13084
rect 19916 13082 19972 13084
rect 19996 13082 20052 13084
rect 19756 13030 19782 13082
rect 19782 13030 19812 13082
rect 19836 13030 19846 13082
rect 19846 13030 19892 13082
rect 19916 13030 19962 13082
rect 19962 13030 19972 13082
rect 19996 13030 20026 13082
rect 20026 13030 20052 13082
rect 19756 13028 19812 13030
rect 19836 13028 19892 13030
rect 19916 13028 19972 13030
rect 19996 13028 20052 13030
rect 18256 11450 18312 11452
rect 18336 11450 18392 11452
rect 18416 11450 18472 11452
rect 18496 11450 18552 11452
rect 18256 11398 18282 11450
rect 18282 11398 18312 11450
rect 18336 11398 18346 11450
rect 18346 11398 18392 11450
rect 18416 11398 18462 11450
rect 18462 11398 18472 11450
rect 18496 11398 18526 11450
rect 18526 11398 18552 11450
rect 18256 11396 18312 11398
rect 18336 11396 18392 11398
rect 18416 11396 18472 11398
rect 18496 11396 18552 11398
rect 19756 11994 19812 11996
rect 19836 11994 19892 11996
rect 19916 11994 19972 11996
rect 19996 11994 20052 11996
rect 19756 11942 19782 11994
rect 19782 11942 19812 11994
rect 19836 11942 19846 11994
rect 19846 11942 19892 11994
rect 19916 11942 19962 11994
rect 19962 11942 19972 11994
rect 19996 11942 20026 11994
rect 20026 11942 20052 11994
rect 19756 11940 19812 11942
rect 19836 11940 19892 11942
rect 19916 11940 19972 11942
rect 19996 11940 20052 11942
rect 18256 10362 18312 10364
rect 18336 10362 18392 10364
rect 18416 10362 18472 10364
rect 18496 10362 18552 10364
rect 18256 10310 18282 10362
rect 18282 10310 18312 10362
rect 18336 10310 18346 10362
rect 18346 10310 18392 10362
rect 18416 10310 18462 10362
rect 18462 10310 18472 10362
rect 18496 10310 18526 10362
rect 18526 10310 18552 10362
rect 18256 10308 18312 10310
rect 18336 10308 18392 10310
rect 18416 10308 18472 10310
rect 18496 10308 18552 10310
rect 18256 9274 18312 9276
rect 18336 9274 18392 9276
rect 18416 9274 18472 9276
rect 18496 9274 18552 9276
rect 18256 9222 18282 9274
rect 18282 9222 18312 9274
rect 18336 9222 18346 9274
rect 18346 9222 18392 9274
rect 18416 9222 18462 9274
rect 18462 9222 18472 9274
rect 18496 9222 18526 9274
rect 18526 9222 18552 9274
rect 18256 9220 18312 9222
rect 18336 9220 18392 9222
rect 18416 9220 18472 9222
rect 18496 9220 18552 9222
rect 16756 8730 16812 8732
rect 16836 8730 16892 8732
rect 16916 8730 16972 8732
rect 16996 8730 17052 8732
rect 16756 8678 16782 8730
rect 16782 8678 16812 8730
rect 16836 8678 16846 8730
rect 16846 8678 16892 8730
rect 16916 8678 16962 8730
rect 16962 8678 16972 8730
rect 16996 8678 17026 8730
rect 17026 8678 17052 8730
rect 16756 8676 16812 8678
rect 16836 8676 16892 8678
rect 16916 8676 16972 8678
rect 16996 8676 17052 8678
rect 16756 7642 16812 7644
rect 16836 7642 16892 7644
rect 16916 7642 16972 7644
rect 16996 7642 17052 7644
rect 16756 7590 16782 7642
rect 16782 7590 16812 7642
rect 16836 7590 16846 7642
rect 16846 7590 16892 7642
rect 16916 7590 16962 7642
rect 16962 7590 16972 7642
rect 16996 7590 17026 7642
rect 17026 7590 17052 7642
rect 16756 7588 16812 7590
rect 16836 7588 16892 7590
rect 16916 7588 16972 7590
rect 16996 7588 17052 7590
rect 16756 6554 16812 6556
rect 16836 6554 16892 6556
rect 16916 6554 16972 6556
rect 16996 6554 17052 6556
rect 16756 6502 16782 6554
rect 16782 6502 16812 6554
rect 16836 6502 16846 6554
rect 16846 6502 16892 6554
rect 16916 6502 16962 6554
rect 16962 6502 16972 6554
rect 16996 6502 17026 6554
rect 17026 6502 17052 6554
rect 16756 6500 16812 6502
rect 16836 6500 16892 6502
rect 16916 6500 16972 6502
rect 16996 6500 17052 6502
rect 16756 5466 16812 5468
rect 16836 5466 16892 5468
rect 16916 5466 16972 5468
rect 16996 5466 17052 5468
rect 16756 5414 16782 5466
rect 16782 5414 16812 5466
rect 16836 5414 16846 5466
rect 16846 5414 16892 5466
rect 16916 5414 16962 5466
rect 16962 5414 16972 5466
rect 16996 5414 17026 5466
rect 17026 5414 17052 5466
rect 16756 5412 16812 5414
rect 16836 5412 16892 5414
rect 16916 5412 16972 5414
rect 16996 5412 17052 5414
rect 16756 4378 16812 4380
rect 16836 4378 16892 4380
rect 16916 4378 16972 4380
rect 16996 4378 17052 4380
rect 16756 4326 16782 4378
rect 16782 4326 16812 4378
rect 16836 4326 16846 4378
rect 16846 4326 16892 4378
rect 16916 4326 16962 4378
rect 16962 4326 16972 4378
rect 16996 4326 17026 4378
rect 17026 4326 17052 4378
rect 16756 4324 16812 4326
rect 16836 4324 16892 4326
rect 16916 4324 16972 4326
rect 16996 4324 17052 4326
rect 18256 8186 18312 8188
rect 18336 8186 18392 8188
rect 18416 8186 18472 8188
rect 18496 8186 18552 8188
rect 18256 8134 18282 8186
rect 18282 8134 18312 8186
rect 18336 8134 18346 8186
rect 18346 8134 18392 8186
rect 18416 8134 18462 8186
rect 18462 8134 18472 8186
rect 18496 8134 18526 8186
rect 18526 8134 18552 8186
rect 18256 8132 18312 8134
rect 18336 8132 18392 8134
rect 18416 8132 18472 8134
rect 18496 8132 18552 8134
rect 18256 7098 18312 7100
rect 18336 7098 18392 7100
rect 18416 7098 18472 7100
rect 18496 7098 18552 7100
rect 18256 7046 18282 7098
rect 18282 7046 18312 7098
rect 18336 7046 18346 7098
rect 18346 7046 18392 7098
rect 18416 7046 18462 7098
rect 18462 7046 18472 7098
rect 18496 7046 18526 7098
rect 18526 7046 18552 7098
rect 18256 7044 18312 7046
rect 18336 7044 18392 7046
rect 18416 7044 18472 7046
rect 18496 7044 18552 7046
rect 18256 6010 18312 6012
rect 18336 6010 18392 6012
rect 18416 6010 18472 6012
rect 18496 6010 18552 6012
rect 18256 5958 18282 6010
rect 18282 5958 18312 6010
rect 18336 5958 18346 6010
rect 18346 5958 18392 6010
rect 18416 5958 18462 6010
rect 18462 5958 18472 6010
rect 18496 5958 18526 6010
rect 18526 5958 18552 6010
rect 18256 5956 18312 5958
rect 18336 5956 18392 5958
rect 18416 5956 18472 5958
rect 18496 5956 18552 5958
rect 18256 4922 18312 4924
rect 18336 4922 18392 4924
rect 18416 4922 18472 4924
rect 18496 4922 18552 4924
rect 18256 4870 18282 4922
rect 18282 4870 18312 4922
rect 18336 4870 18346 4922
rect 18346 4870 18392 4922
rect 18416 4870 18462 4922
rect 18462 4870 18472 4922
rect 18496 4870 18526 4922
rect 18526 4870 18552 4922
rect 18256 4868 18312 4870
rect 18336 4868 18392 4870
rect 18416 4868 18472 4870
rect 18496 4868 18552 4870
rect 19756 10906 19812 10908
rect 19836 10906 19892 10908
rect 19916 10906 19972 10908
rect 19996 10906 20052 10908
rect 19756 10854 19782 10906
rect 19782 10854 19812 10906
rect 19836 10854 19846 10906
rect 19846 10854 19892 10906
rect 19916 10854 19962 10906
rect 19962 10854 19972 10906
rect 19996 10854 20026 10906
rect 20026 10854 20052 10906
rect 19756 10852 19812 10854
rect 19836 10852 19892 10854
rect 19916 10852 19972 10854
rect 19996 10852 20052 10854
rect 19756 9818 19812 9820
rect 19836 9818 19892 9820
rect 19916 9818 19972 9820
rect 19996 9818 20052 9820
rect 19756 9766 19782 9818
rect 19782 9766 19812 9818
rect 19836 9766 19846 9818
rect 19846 9766 19892 9818
rect 19916 9766 19962 9818
rect 19962 9766 19972 9818
rect 19996 9766 20026 9818
rect 20026 9766 20052 9818
rect 19756 9764 19812 9766
rect 19836 9764 19892 9766
rect 19916 9764 19972 9766
rect 19996 9764 20052 9766
rect 22756 15258 22812 15260
rect 22836 15258 22892 15260
rect 22916 15258 22972 15260
rect 22996 15258 23052 15260
rect 22756 15206 22782 15258
rect 22782 15206 22812 15258
rect 22836 15206 22846 15258
rect 22846 15206 22892 15258
rect 22916 15206 22962 15258
rect 22962 15206 22972 15258
rect 22996 15206 23026 15258
rect 23026 15206 23052 15258
rect 22756 15204 22812 15206
rect 22836 15204 22892 15206
rect 22916 15204 22972 15206
rect 22996 15204 23052 15206
rect 21256 14714 21312 14716
rect 21336 14714 21392 14716
rect 21416 14714 21472 14716
rect 21496 14714 21552 14716
rect 21256 14662 21282 14714
rect 21282 14662 21312 14714
rect 21336 14662 21346 14714
rect 21346 14662 21392 14714
rect 21416 14662 21462 14714
rect 21462 14662 21472 14714
rect 21496 14662 21526 14714
rect 21526 14662 21552 14714
rect 21256 14660 21312 14662
rect 21336 14660 21392 14662
rect 21416 14660 21472 14662
rect 21496 14660 21552 14662
rect 21638 14456 21694 14512
rect 25756 27226 25812 27228
rect 25836 27226 25892 27228
rect 25916 27226 25972 27228
rect 25996 27226 26052 27228
rect 25756 27174 25782 27226
rect 25782 27174 25812 27226
rect 25836 27174 25846 27226
rect 25846 27174 25892 27226
rect 25916 27174 25962 27226
rect 25962 27174 25972 27226
rect 25996 27174 26026 27226
rect 26026 27174 26052 27226
rect 25756 27172 25812 27174
rect 25836 27172 25892 27174
rect 25916 27172 25972 27174
rect 25996 27172 26052 27174
rect 24256 26682 24312 26684
rect 24336 26682 24392 26684
rect 24416 26682 24472 26684
rect 24496 26682 24552 26684
rect 24256 26630 24282 26682
rect 24282 26630 24312 26682
rect 24336 26630 24346 26682
rect 24346 26630 24392 26682
rect 24416 26630 24462 26682
rect 24462 26630 24472 26682
rect 24496 26630 24526 26682
rect 24526 26630 24552 26682
rect 24256 26628 24312 26630
rect 24336 26628 24392 26630
rect 24416 26628 24472 26630
rect 24496 26628 24552 26630
rect 27256 26682 27312 26684
rect 27336 26682 27392 26684
rect 27416 26682 27472 26684
rect 27496 26682 27552 26684
rect 27256 26630 27282 26682
rect 27282 26630 27312 26682
rect 27336 26630 27346 26682
rect 27346 26630 27392 26682
rect 27416 26630 27462 26682
rect 27462 26630 27472 26682
rect 27496 26630 27526 26682
rect 27526 26630 27552 26682
rect 27256 26628 27312 26630
rect 27336 26628 27392 26630
rect 27416 26628 27472 26630
rect 27496 26628 27552 26630
rect 25756 26138 25812 26140
rect 25836 26138 25892 26140
rect 25916 26138 25972 26140
rect 25996 26138 26052 26140
rect 25756 26086 25782 26138
rect 25782 26086 25812 26138
rect 25836 26086 25846 26138
rect 25846 26086 25892 26138
rect 25916 26086 25962 26138
rect 25962 26086 25972 26138
rect 25996 26086 26026 26138
rect 26026 26086 26052 26138
rect 25756 26084 25812 26086
rect 25836 26084 25892 26086
rect 25916 26084 25972 26086
rect 25996 26084 26052 26086
rect 24256 25594 24312 25596
rect 24336 25594 24392 25596
rect 24416 25594 24472 25596
rect 24496 25594 24552 25596
rect 24256 25542 24282 25594
rect 24282 25542 24312 25594
rect 24336 25542 24346 25594
rect 24346 25542 24392 25594
rect 24416 25542 24462 25594
rect 24462 25542 24472 25594
rect 24496 25542 24526 25594
rect 24526 25542 24552 25594
rect 24256 25540 24312 25542
rect 24336 25540 24392 25542
rect 24416 25540 24472 25542
rect 24496 25540 24552 25542
rect 27256 25594 27312 25596
rect 27336 25594 27392 25596
rect 27416 25594 27472 25596
rect 27496 25594 27552 25596
rect 27256 25542 27282 25594
rect 27282 25542 27312 25594
rect 27336 25542 27346 25594
rect 27346 25542 27392 25594
rect 27416 25542 27462 25594
rect 27462 25542 27472 25594
rect 27496 25542 27526 25594
rect 27526 25542 27552 25594
rect 27256 25540 27312 25542
rect 27336 25540 27392 25542
rect 27416 25540 27472 25542
rect 27496 25540 27552 25542
rect 25756 25050 25812 25052
rect 25836 25050 25892 25052
rect 25916 25050 25972 25052
rect 25996 25050 26052 25052
rect 25756 24998 25782 25050
rect 25782 24998 25812 25050
rect 25836 24998 25846 25050
rect 25846 24998 25892 25050
rect 25916 24998 25962 25050
rect 25962 24998 25972 25050
rect 25996 24998 26026 25050
rect 26026 24998 26052 25050
rect 25756 24996 25812 24998
rect 25836 24996 25892 24998
rect 25916 24996 25972 24998
rect 25996 24996 26052 24998
rect 24256 24506 24312 24508
rect 24336 24506 24392 24508
rect 24416 24506 24472 24508
rect 24496 24506 24552 24508
rect 24256 24454 24282 24506
rect 24282 24454 24312 24506
rect 24336 24454 24346 24506
rect 24346 24454 24392 24506
rect 24416 24454 24462 24506
rect 24462 24454 24472 24506
rect 24496 24454 24526 24506
rect 24526 24454 24552 24506
rect 24256 24452 24312 24454
rect 24336 24452 24392 24454
rect 24416 24452 24472 24454
rect 24496 24452 24552 24454
rect 27256 24506 27312 24508
rect 27336 24506 27392 24508
rect 27416 24506 27472 24508
rect 27496 24506 27552 24508
rect 27256 24454 27282 24506
rect 27282 24454 27312 24506
rect 27336 24454 27346 24506
rect 27346 24454 27392 24506
rect 27416 24454 27462 24506
rect 27462 24454 27472 24506
rect 27496 24454 27526 24506
rect 27526 24454 27552 24506
rect 27256 24452 27312 24454
rect 27336 24452 27392 24454
rect 27416 24452 27472 24454
rect 27496 24452 27552 24454
rect 25756 23962 25812 23964
rect 25836 23962 25892 23964
rect 25916 23962 25972 23964
rect 25996 23962 26052 23964
rect 25756 23910 25782 23962
rect 25782 23910 25812 23962
rect 25836 23910 25846 23962
rect 25846 23910 25892 23962
rect 25916 23910 25962 23962
rect 25962 23910 25972 23962
rect 25996 23910 26026 23962
rect 26026 23910 26052 23962
rect 25756 23908 25812 23910
rect 25836 23908 25892 23910
rect 25916 23908 25972 23910
rect 25996 23908 26052 23910
rect 24256 23418 24312 23420
rect 24336 23418 24392 23420
rect 24416 23418 24472 23420
rect 24496 23418 24552 23420
rect 24256 23366 24282 23418
rect 24282 23366 24312 23418
rect 24336 23366 24346 23418
rect 24346 23366 24392 23418
rect 24416 23366 24462 23418
rect 24462 23366 24472 23418
rect 24496 23366 24526 23418
rect 24526 23366 24552 23418
rect 24256 23364 24312 23366
rect 24336 23364 24392 23366
rect 24416 23364 24472 23366
rect 24496 23364 24552 23366
rect 27256 23418 27312 23420
rect 27336 23418 27392 23420
rect 27416 23418 27472 23420
rect 27496 23418 27552 23420
rect 27256 23366 27282 23418
rect 27282 23366 27312 23418
rect 27336 23366 27346 23418
rect 27346 23366 27392 23418
rect 27416 23366 27462 23418
rect 27462 23366 27472 23418
rect 27496 23366 27526 23418
rect 27526 23366 27552 23418
rect 27256 23364 27312 23366
rect 27336 23364 27392 23366
rect 27416 23364 27472 23366
rect 27496 23364 27552 23366
rect 25756 22874 25812 22876
rect 25836 22874 25892 22876
rect 25916 22874 25972 22876
rect 25996 22874 26052 22876
rect 25756 22822 25782 22874
rect 25782 22822 25812 22874
rect 25836 22822 25846 22874
rect 25846 22822 25892 22874
rect 25916 22822 25962 22874
rect 25962 22822 25972 22874
rect 25996 22822 26026 22874
rect 26026 22822 26052 22874
rect 25756 22820 25812 22822
rect 25836 22820 25892 22822
rect 25916 22820 25972 22822
rect 25996 22820 26052 22822
rect 24256 22330 24312 22332
rect 24336 22330 24392 22332
rect 24416 22330 24472 22332
rect 24496 22330 24552 22332
rect 24256 22278 24282 22330
rect 24282 22278 24312 22330
rect 24336 22278 24346 22330
rect 24346 22278 24392 22330
rect 24416 22278 24462 22330
rect 24462 22278 24472 22330
rect 24496 22278 24526 22330
rect 24526 22278 24552 22330
rect 24256 22276 24312 22278
rect 24336 22276 24392 22278
rect 24416 22276 24472 22278
rect 24496 22276 24552 22278
rect 27256 22330 27312 22332
rect 27336 22330 27392 22332
rect 27416 22330 27472 22332
rect 27496 22330 27552 22332
rect 27256 22278 27282 22330
rect 27282 22278 27312 22330
rect 27336 22278 27346 22330
rect 27346 22278 27392 22330
rect 27416 22278 27462 22330
rect 27462 22278 27472 22330
rect 27496 22278 27526 22330
rect 27526 22278 27552 22330
rect 27256 22276 27312 22278
rect 27336 22276 27392 22278
rect 27416 22276 27472 22278
rect 27496 22276 27552 22278
rect 25756 21786 25812 21788
rect 25836 21786 25892 21788
rect 25916 21786 25972 21788
rect 25996 21786 26052 21788
rect 25756 21734 25782 21786
rect 25782 21734 25812 21786
rect 25836 21734 25846 21786
rect 25846 21734 25892 21786
rect 25916 21734 25962 21786
rect 25962 21734 25972 21786
rect 25996 21734 26026 21786
rect 26026 21734 26052 21786
rect 25756 21732 25812 21734
rect 25836 21732 25892 21734
rect 25916 21732 25972 21734
rect 25996 21732 26052 21734
rect 24256 21242 24312 21244
rect 24336 21242 24392 21244
rect 24416 21242 24472 21244
rect 24496 21242 24552 21244
rect 24256 21190 24282 21242
rect 24282 21190 24312 21242
rect 24336 21190 24346 21242
rect 24346 21190 24392 21242
rect 24416 21190 24462 21242
rect 24462 21190 24472 21242
rect 24496 21190 24526 21242
rect 24526 21190 24552 21242
rect 24256 21188 24312 21190
rect 24336 21188 24392 21190
rect 24416 21188 24472 21190
rect 24496 21188 24552 21190
rect 27256 21242 27312 21244
rect 27336 21242 27392 21244
rect 27416 21242 27472 21244
rect 27496 21242 27552 21244
rect 27256 21190 27282 21242
rect 27282 21190 27312 21242
rect 27336 21190 27346 21242
rect 27346 21190 27392 21242
rect 27416 21190 27462 21242
rect 27462 21190 27472 21242
rect 27496 21190 27526 21242
rect 27526 21190 27552 21242
rect 27256 21188 27312 21190
rect 27336 21188 27392 21190
rect 27416 21188 27472 21190
rect 27496 21188 27552 21190
rect 25756 20698 25812 20700
rect 25836 20698 25892 20700
rect 25916 20698 25972 20700
rect 25996 20698 26052 20700
rect 25756 20646 25782 20698
rect 25782 20646 25812 20698
rect 25836 20646 25846 20698
rect 25846 20646 25892 20698
rect 25916 20646 25962 20698
rect 25962 20646 25972 20698
rect 25996 20646 26026 20698
rect 26026 20646 26052 20698
rect 25756 20644 25812 20646
rect 25836 20644 25892 20646
rect 25916 20644 25972 20646
rect 25996 20644 26052 20646
rect 24256 20154 24312 20156
rect 24336 20154 24392 20156
rect 24416 20154 24472 20156
rect 24496 20154 24552 20156
rect 24256 20102 24282 20154
rect 24282 20102 24312 20154
rect 24336 20102 24346 20154
rect 24346 20102 24392 20154
rect 24416 20102 24462 20154
rect 24462 20102 24472 20154
rect 24496 20102 24526 20154
rect 24526 20102 24552 20154
rect 24256 20100 24312 20102
rect 24336 20100 24392 20102
rect 24416 20100 24472 20102
rect 24496 20100 24552 20102
rect 27256 20154 27312 20156
rect 27336 20154 27392 20156
rect 27416 20154 27472 20156
rect 27496 20154 27552 20156
rect 27256 20102 27282 20154
rect 27282 20102 27312 20154
rect 27336 20102 27346 20154
rect 27346 20102 27392 20154
rect 27416 20102 27462 20154
rect 27462 20102 27472 20154
rect 27496 20102 27526 20154
rect 27526 20102 27552 20154
rect 27256 20100 27312 20102
rect 27336 20100 27392 20102
rect 27416 20100 27472 20102
rect 27496 20100 27552 20102
rect 25756 19610 25812 19612
rect 25836 19610 25892 19612
rect 25916 19610 25972 19612
rect 25996 19610 26052 19612
rect 25756 19558 25782 19610
rect 25782 19558 25812 19610
rect 25836 19558 25846 19610
rect 25846 19558 25892 19610
rect 25916 19558 25962 19610
rect 25962 19558 25972 19610
rect 25996 19558 26026 19610
rect 26026 19558 26052 19610
rect 25756 19556 25812 19558
rect 25836 19556 25892 19558
rect 25916 19556 25972 19558
rect 25996 19556 26052 19558
rect 24256 19066 24312 19068
rect 24336 19066 24392 19068
rect 24416 19066 24472 19068
rect 24496 19066 24552 19068
rect 24256 19014 24282 19066
rect 24282 19014 24312 19066
rect 24336 19014 24346 19066
rect 24346 19014 24392 19066
rect 24416 19014 24462 19066
rect 24462 19014 24472 19066
rect 24496 19014 24526 19066
rect 24526 19014 24552 19066
rect 24256 19012 24312 19014
rect 24336 19012 24392 19014
rect 24416 19012 24472 19014
rect 24496 19012 24552 19014
rect 27256 19066 27312 19068
rect 27336 19066 27392 19068
rect 27416 19066 27472 19068
rect 27496 19066 27552 19068
rect 27256 19014 27282 19066
rect 27282 19014 27312 19066
rect 27336 19014 27346 19066
rect 27346 19014 27392 19066
rect 27416 19014 27462 19066
rect 27462 19014 27472 19066
rect 27496 19014 27526 19066
rect 27526 19014 27552 19066
rect 27256 19012 27312 19014
rect 27336 19012 27392 19014
rect 27416 19012 27472 19014
rect 27496 19012 27552 19014
rect 25756 18522 25812 18524
rect 25836 18522 25892 18524
rect 25916 18522 25972 18524
rect 25996 18522 26052 18524
rect 25756 18470 25782 18522
rect 25782 18470 25812 18522
rect 25836 18470 25846 18522
rect 25846 18470 25892 18522
rect 25916 18470 25962 18522
rect 25962 18470 25972 18522
rect 25996 18470 26026 18522
rect 26026 18470 26052 18522
rect 25756 18468 25812 18470
rect 25836 18468 25892 18470
rect 25916 18468 25972 18470
rect 25996 18468 26052 18470
rect 24256 17978 24312 17980
rect 24336 17978 24392 17980
rect 24416 17978 24472 17980
rect 24496 17978 24552 17980
rect 24256 17926 24282 17978
rect 24282 17926 24312 17978
rect 24336 17926 24346 17978
rect 24346 17926 24392 17978
rect 24416 17926 24462 17978
rect 24462 17926 24472 17978
rect 24496 17926 24526 17978
rect 24526 17926 24552 17978
rect 24256 17924 24312 17926
rect 24336 17924 24392 17926
rect 24416 17924 24472 17926
rect 24496 17924 24552 17926
rect 27256 17978 27312 17980
rect 27336 17978 27392 17980
rect 27416 17978 27472 17980
rect 27496 17978 27552 17980
rect 27256 17926 27282 17978
rect 27282 17926 27312 17978
rect 27336 17926 27346 17978
rect 27346 17926 27392 17978
rect 27416 17926 27462 17978
rect 27462 17926 27472 17978
rect 27496 17926 27526 17978
rect 27526 17926 27552 17978
rect 27256 17924 27312 17926
rect 27336 17924 27392 17926
rect 27416 17924 27472 17926
rect 27496 17924 27552 17926
rect 25756 17434 25812 17436
rect 25836 17434 25892 17436
rect 25916 17434 25972 17436
rect 25996 17434 26052 17436
rect 25756 17382 25782 17434
rect 25782 17382 25812 17434
rect 25836 17382 25846 17434
rect 25846 17382 25892 17434
rect 25916 17382 25962 17434
rect 25962 17382 25972 17434
rect 25996 17382 26026 17434
rect 26026 17382 26052 17434
rect 25756 17380 25812 17382
rect 25836 17380 25892 17382
rect 25916 17380 25972 17382
rect 25996 17380 26052 17382
rect 24256 16890 24312 16892
rect 24336 16890 24392 16892
rect 24416 16890 24472 16892
rect 24496 16890 24552 16892
rect 24256 16838 24282 16890
rect 24282 16838 24312 16890
rect 24336 16838 24346 16890
rect 24346 16838 24392 16890
rect 24416 16838 24462 16890
rect 24462 16838 24472 16890
rect 24496 16838 24526 16890
rect 24526 16838 24552 16890
rect 24256 16836 24312 16838
rect 24336 16836 24392 16838
rect 24416 16836 24472 16838
rect 24496 16836 24552 16838
rect 27256 16890 27312 16892
rect 27336 16890 27392 16892
rect 27416 16890 27472 16892
rect 27496 16890 27552 16892
rect 27256 16838 27282 16890
rect 27282 16838 27312 16890
rect 27336 16838 27346 16890
rect 27346 16838 27392 16890
rect 27416 16838 27462 16890
rect 27462 16838 27472 16890
rect 27496 16838 27526 16890
rect 27526 16838 27552 16890
rect 27256 16836 27312 16838
rect 27336 16836 27392 16838
rect 27416 16836 27472 16838
rect 27496 16836 27552 16838
rect 25756 16346 25812 16348
rect 25836 16346 25892 16348
rect 25916 16346 25972 16348
rect 25996 16346 26052 16348
rect 25756 16294 25782 16346
rect 25782 16294 25812 16346
rect 25836 16294 25846 16346
rect 25846 16294 25892 16346
rect 25916 16294 25962 16346
rect 25962 16294 25972 16346
rect 25996 16294 26026 16346
rect 26026 16294 26052 16346
rect 25756 16292 25812 16294
rect 25836 16292 25892 16294
rect 25916 16292 25972 16294
rect 25996 16292 26052 16294
rect 24256 15802 24312 15804
rect 24336 15802 24392 15804
rect 24416 15802 24472 15804
rect 24496 15802 24552 15804
rect 24256 15750 24282 15802
rect 24282 15750 24312 15802
rect 24336 15750 24346 15802
rect 24346 15750 24392 15802
rect 24416 15750 24462 15802
rect 24462 15750 24472 15802
rect 24496 15750 24526 15802
rect 24526 15750 24552 15802
rect 24256 15748 24312 15750
rect 24336 15748 24392 15750
rect 24416 15748 24472 15750
rect 24496 15748 24552 15750
rect 27256 15802 27312 15804
rect 27336 15802 27392 15804
rect 27416 15802 27472 15804
rect 27496 15802 27552 15804
rect 27256 15750 27282 15802
rect 27282 15750 27312 15802
rect 27336 15750 27346 15802
rect 27346 15750 27392 15802
rect 27416 15750 27462 15802
rect 27462 15750 27472 15802
rect 27496 15750 27526 15802
rect 27526 15750 27552 15802
rect 27256 15748 27312 15750
rect 27336 15748 27392 15750
rect 27416 15748 27472 15750
rect 27496 15748 27552 15750
rect 25756 15258 25812 15260
rect 25836 15258 25892 15260
rect 25916 15258 25972 15260
rect 25996 15258 26052 15260
rect 25756 15206 25782 15258
rect 25782 15206 25812 15258
rect 25836 15206 25846 15258
rect 25846 15206 25892 15258
rect 25916 15206 25962 15258
rect 25962 15206 25972 15258
rect 25996 15206 26026 15258
rect 26026 15206 26052 15258
rect 25756 15204 25812 15206
rect 25836 15204 25892 15206
rect 25916 15204 25972 15206
rect 25996 15204 26052 15206
rect 24256 14714 24312 14716
rect 24336 14714 24392 14716
rect 24416 14714 24472 14716
rect 24496 14714 24552 14716
rect 24256 14662 24282 14714
rect 24282 14662 24312 14714
rect 24336 14662 24346 14714
rect 24346 14662 24392 14714
rect 24416 14662 24462 14714
rect 24462 14662 24472 14714
rect 24496 14662 24526 14714
rect 24526 14662 24552 14714
rect 24256 14660 24312 14662
rect 24336 14660 24392 14662
rect 24416 14660 24472 14662
rect 24496 14660 24552 14662
rect 27256 14714 27312 14716
rect 27336 14714 27392 14716
rect 27416 14714 27472 14716
rect 27496 14714 27552 14716
rect 27256 14662 27282 14714
rect 27282 14662 27312 14714
rect 27336 14662 27346 14714
rect 27346 14662 27392 14714
rect 27416 14662 27462 14714
rect 27462 14662 27472 14714
rect 27496 14662 27526 14714
rect 27526 14662 27552 14714
rect 27256 14660 27312 14662
rect 27336 14660 27392 14662
rect 27416 14660 27472 14662
rect 27496 14660 27552 14662
rect 21256 13626 21312 13628
rect 21336 13626 21392 13628
rect 21416 13626 21472 13628
rect 21496 13626 21552 13628
rect 21256 13574 21282 13626
rect 21282 13574 21312 13626
rect 21336 13574 21346 13626
rect 21346 13574 21392 13626
rect 21416 13574 21462 13626
rect 21462 13574 21472 13626
rect 21496 13574 21526 13626
rect 21526 13574 21552 13626
rect 21256 13572 21312 13574
rect 21336 13572 21392 13574
rect 21416 13572 21472 13574
rect 21496 13572 21552 13574
rect 21256 12538 21312 12540
rect 21336 12538 21392 12540
rect 21416 12538 21472 12540
rect 21496 12538 21552 12540
rect 21256 12486 21282 12538
rect 21282 12486 21312 12538
rect 21336 12486 21346 12538
rect 21346 12486 21392 12538
rect 21416 12486 21462 12538
rect 21462 12486 21472 12538
rect 21496 12486 21526 12538
rect 21526 12486 21552 12538
rect 21256 12484 21312 12486
rect 21336 12484 21392 12486
rect 21416 12484 21472 12486
rect 21496 12484 21552 12486
rect 21256 11450 21312 11452
rect 21336 11450 21392 11452
rect 21416 11450 21472 11452
rect 21496 11450 21552 11452
rect 21256 11398 21282 11450
rect 21282 11398 21312 11450
rect 21336 11398 21346 11450
rect 21346 11398 21392 11450
rect 21416 11398 21462 11450
rect 21462 11398 21472 11450
rect 21496 11398 21526 11450
rect 21526 11398 21552 11450
rect 21256 11396 21312 11398
rect 21336 11396 21392 11398
rect 21416 11396 21472 11398
rect 21496 11396 21552 11398
rect 21256 10362 21312 10364
rect 21336 10362 21392 10364
rect 21416 10362 21472 10364
rect 21496 10362 21552 10364
rect 21256 10310 21282 10362
rect 21282 10310 21312 10362
rect 21336 10310 21346 10362
rect 21346 10310 21392 10362
rect 21416 10310 21462 10362
rect 21462 10310 21472 10362
rect 21496 10310 21526 10362
rect 21526 10310 21552 10362
rect 21256 10308 21312 10310
rect 21336 10308 21392 10310
rect 21416 10308 21472 10310
rect 21496 10308 21552 10310
rect 20994 9968 21050 10024
rect 19756 8730 19812 8732
rect 19836 8730 19892 8732
rect 19916 8730 19972 8732
rect 19996 8730 20052 8732
rect 19756 8678 19782 8730
rect 19782 8678 19812 8730
rect 19836 8678 19846 8730
rect 19846 8678 19892 8730
rect 19916 8678 19962 8730
rect 19962 8678 19972 8730
rect 19996 8678 20026 8730
rect 20026 8678 20052 8730
rect 19756 8676 19812 8678
rect 19836 8676 19892 8678
rect 19916 8676 19972 8678
rect 19996 8676 20052 8678
rect 21256 9274 21312 9276
rect 21336 9274 21392 9276
rect 21416 9274 21472 9276
rect 21496 9274 21552 9276
rect 21256 9222 21282 9274
rect 21282 9222 21312 9274
rect 21336 9222 21346 9274
rect 21346 9222 21392 9274
rect 21416 9222 21462 9274
rect 21462 9222 21472 9274
rect 21496 9222 21526 9274
rect 21526 9222 21552 9274
rect 21256 9220 21312 9222
rect 21336 9220 21392 9222
rect 21416 9220 21472 9222
rect 21496 9220 21552 9222
rect 22756 14170 22812 14172
rect 22836 14170 22892 14172
rect 22916 14170 22972 14172
rect 22996 14170 23052 14172
rect 22756 14118 22782 14170
rect 22782 14118 22812 14170
rect 22836 14118 22846 14170
rect 22846 14118 22892 14170
rect 22916 14118 22962 14170
rect 22962 14118 22972 14170
rect 22996 14118 23026 14170
rect 23026 14118 23052 14170
rect 22756 14116 22812 14118
rect 22836 14116 22892 14118
rect 22916 14116 22972 14118
rect 22996 14116 23052 14118
rect 25756 14170 25812 14172
rect 25836 14170 25892 14172
rect 25916 14170 25972 14172
rect 25996 14170 26052 14172
rect 25756 14118 25782 14170
rect 25782 14118 25812 14170
rect 25836 14118 25846 14170
rect 25846 14118 25892 14170
rect 25916 14118 25962 14170
rect 25962 14118 25972 14170
rect 25996 14118 26026 14170
rect 26026 14118 26052 14170
rect 25756 14116 25812 14118
rect 25836 14116 25892 14118
rect 25916 14116 25972 14118
rect 25996 14116 26052 14118
rect 24256 13626 24312 13628
rect 24336 13626 24392 13628
rect 24416 13626 24472 13628
rect 24496 13626 24552 13628
rect 24256 13574 24282 13626
rect 24282 13574 24312 13626
rect 24336 13574 24346 13626
rect 24346 13574 24392 13626
rect 24416 13574 24462 13626
rect 24462 13574 24472 13626
rect 24496 13574 24526 13626
rect 24526 13574 24552 13626
rect 24256 13572 24312 13574
rect 24336 13572 24392 13574
rect 24416 13572 24472 13574
rect 24496 13572 24552 13574
rect 27256 13626 27312 13628
rect 27336 13626 27392 13628
rect 27416 13626 27472 13628
rect 27496 13626 27552 13628
rect 27256 13574 27282 13626
rect 27282 13574 27312 13626
rect 27336 13574 27346 13626
rect 27346 13574 27392 13626
rect 27416 13574 27462 13626
rect 27462 13574 27472 13626
rect 27496 13574 27526 13626
rect 27526 13574 27552 13626
rect 27256 13572 27312 13574
rect 27336 13572 27392 13574
rect 27416 13572 27472 13574
rect 27496 13572 27552 13574
rect 22756 13082 22812 13084
rect 22836 13082 22892 13084
rect 22916 13082 22972 13084
rect 22996 13082 23052 13084
rect 22756 13030 22782 13082
rect 22782 13030 22812 13082
rect 22836 13030 22846 13082
rect 22846 13030 22892 13082
rect 22916 13030 22962 13082
rect 22962 13030 22972 13082
rect 22996 13030 23026 13082
rect 23026 13030 23052 13082
rect 22756 13028 22812 13030
rect 22836 13028 22892 13030
rect 22916 13028 22972 13030
rect 22996 13028 23052 13030
rect 23202 12688 23258 12744
rect 25756 13082 25812 13084
rect 25836 13082 25892 13084
rect 25916 13082 25972 13084
rect 25996 13082 26052 13084
rect 25756 13030 25782 13082
rect 25782 13030 25812 13082
rect 25836 13030 25846 13082
rect 25846 13030 25892 13082
rect 25916 13030 25962 13082
rect 25962 13030 25972 13082
rect 25996 13030 26026 13082
rect 26026 13030 26052 13082
rect 25756 13028 25812 13030
rect 25836 13028 25892 13030
rect 25916 13028 25972 13030
rect 25996 13028 26052 13030
rect 24256 12538 24312 12540
rect 24336 12538 24392 12540
rect 24416 12538 24472 12540
rect 24496 12538 24552 12540
rect 24256 12486 24282 12538
rect 24282 12486 24312 12538
rect 24336 12486 24346 12538
rect 24346 12486 24392 12538
rect 24416 12486 24462 12538
rect 24462 12486 24472 12538
rect 24496 12486 24526 12538
rect 24526 12486 24552 12538
rect 24256 12484 24312 12486
rect 24336 12484 24392 12486
rect 24416 12484 24472 12486
rect 24496 12484 24552 12486
rect 27256 12538 27312 12540
rect 27336 12538 27392 12540
rect 27416 12538 27472 12540
rect 27496 12538 27552 12540
rect 27256 12486 27282 12538
rect 27282 12486 27312 12538
rect 27336 12486 27346 12538
rect 27346 12486 27392 12538
rect 27416 12486 27462 12538
rect 27462 12486 27472 12538
rect 27496 12486 27526 12538
rect 27526 12486 27552 12538
rect 27256 12484 27312 12486
rect 27336 12484 27392 12486
rect 27416 12484 27472 12486
rect 27496 12484 27552 12486
rect 22756 11994 22812 11996
rect 22836 11994 22892 11996
rect 22916 11994 22972 11996
rect 22996 11994 23052 11996
rect 22756 11942 22782 11994
rect 22782 11942 22812 11994
rect 22836 11942 22846 11994
rect 22846 11942 22892 11994
rect 22916 11942 22962 11994
rect 22962 11942 22972 11994
rect 22996 11942 23026 11994
rect 23026 11942 23052 11994
rect 22756 11940 22812 11942
rect 22836 11940 22892 11942
rect 22916 11940 22972 11942
rect 22996 11940 23052 11942
rect 25756 11994 25812 11996
rect 25836 11994 25892 11996
rect 25916 11994 25972 11996
rect 25996 11994 26052 11996
rect 25756 11942 25782 11994
rect 25782 11942 25812 11994
rect 25836 11942 25846 11994
rect 25846 11942 25892 11994
rect 25916 11942 25962 11994
rect 25962 11942 25972 11994
rect 25996 11942 26026 11994
rect 26026 11942 26052 11994
rect 25756 11940 25812 11942
rect 25836 11940 25892 11942
rect 25916 11940 25972 11942
rect 25996 11940 26052 11942
rect 24256 11450 24312 11452
rect 24336 11450 24392 11452
rect 24416 11450 24472 11452
rect 24496 11450 24552 11452
rect 24256 11398 24282 11450
rect 24282 11398 24312 11450
rect 24336 11398 24346 11450
rect 24346 11398 24392 11450
rect 24416 11398 24462 11450
rect 24462 11398 24472 11450
rect 24496 11398 24526 11450
rect 24526 11398 24552 11450
rect 24256 11396 24312 11398
rect 24336 11396 24392 11398
rect 24416 11396 24472 11398
rect 24496 11396 24552 11398
rect 27256 11450 27312 11452
rect 27336 11450 27392 11452
rect 27416 11450 27472 11452
rect 27496 11450 27552 11452
rect 27256 11398 27282 11450
rect 27282 11398 27312 11450
rect 27336 11398 27346 11450
rect 27346 11398 27392 11450
rect 27416 11398 27462 11450
rect 27462 11398 27472 11450
rect 27496 11398 27526 11450
rect 27526 11398 27552 11450
rect 27256 11396 27312 11398
rect 27336 11396 27392 11398
rect 27416 11396 27472 11398
rect 27496 11396 27552 11398
rect 28722 11056 28778 11112
rect 22756 10906 22812 10908
rect 22836 10906 22892 10908
rect 22916 10906 22972 10908
rect 22996 10906 23052 10908
rect 22756 10854 22782 10906
rect 22782 10854 22812 10906
rect 22836 10854 22846 10906
rect 22846 10854 22892 10906
rect 22916 10854 22962 10906
rect 22962 10854 22972 10906
rect 22996 10854 23026 10906
rect 23026 10854 23052 10906
rect 22756 10852 22812 10854
rect 22836 10852 22892 10854
rect 22916 10852 22972 10854
rect 22996 10852 23052 10854
rect 25756 10906 25812 10908
rect 25836 10906 25892 10908
rect 25916 10906 25972 10908
rect 25996 10906 26052 10908
rect 25756 10854 25782 10906
rect 25782 10854 25812 10906
rect 25836 10854 25846 10906
rect 25846 10854 25892 10906
rect 25916 10854 25962 10906
rect 25962 10854 25972 10906
rect 25996 10854 26026 10906
rect 26026 10854 26052 10906
rect 25756 10852 25812 10854
rect 25836 10852 25892 10854
rect 25916 10852 25972 10854
rect 25996 10852 26052 10854
rect 19756 7642 19812 7644
rect 19836 7642 19892 7644
rect 19916 7642 19972 7644
rect 19996 7642 20052 7644
rect 19756 7590 19782 7642
rect 19782 7590 19812 7642
rect 19836 7590 19846 7642
rect 19846 7590 19892 7642
rect 19916 7590 19962 7642
rect 19962 7590 19972 7642
rect 19996 7590 20026 7642
rect 20026 7590 20052 7642
rect 19756 7588 19812 7590
rect 19836 7588 19892 7590
rect 19916 7588 19972 7590
rect 19996 7588 20052 7590
rect 19756 6554 19812 6556
rect 19836 6554 19892 6556
rect 19916 6554 19972 6556
rect 19996 6554 20052 6556
rect 19756 6502 19782 6554
rect 19782 6502 19812 6554
rect 19836 6502 19846 6554
rect 19846 6502 19892 6554
rect 19916 6502 19962 6554
rect 19962 6502 19972 6554
rect 19996 6502 20026 6554
rect 20026 6502 20052 6554
rect 19756 6500 19812 6502
rect 19836 6500 19892 6502
rect 19916 6500 19972 6502
rect 19996 6500 20052 6502
rect 19756 5466 19812 5468
rect 19836 5466 19892 5468
rect 19916 5466 19972 5468
rect 19996 5466 20052 5468
rect 19756 5414 19782 5466
rect 19782 5414 19812 5466
rect 19836 5414 19846 5466
rect 19846 5414 19892 5466
rect 19916 5414 19962 5466
rect 19962 5414 19972 5466
rect 19996 5414 20026 5466
rect 20026 5414 20052 5466
rect 19756 5412 19812 5414
rect 19836 5412 19892 5414
rect 19916 5412 19972 5414
rect 19996 5412 20052 5414
rect 21256 8186 21312 8188
rect 21336 8186 21392 8188
rect 21416 8186 21472 8188
rect 21496 8186 21552 8188
rect 21256 8134 21282 8186
rect 21282 8134 21312 8186
rect 21336 8134 21346 8186
rect 21346 8134 21392 8186
rect 21416 8134 21462 8186
rect 21462 8134 21472 8186
rect 21496 8134 21526 8186
rect 21526 8134 21552 8186
rect 21256 8132 21312 8134
rect 21336 8132 21392 8134
rect 21416 8132 21472 8134
rect 21496 8132 21552 8134
rect 21256 7098 21312 7100
rect 21336 7098 21392 7100
rect 21416 7098 21472 7100
rect 21496 7098 21552 7100
rect 21256 7046 21282 7098
rect 21282 7046 21312 7098
rect 21336 7046 21346 7098
rect 21346 7046 21392 7098
rect 21416 7046 21462 7098
rect 21462 7046 21472 7098
rect 21496 7046 21526 7098
rect 21526 7046 21552 7098
rect 21256 7044 21312 7046
rect 21336 7044 21392 7046
rect 21416 7044 21472 7046
rect 21496 7044 21552 7046
rect 24256 10362 24312 10364
rect 24336 10362 24392 10364
rect 24416 10362 24472 10364
rect 24496 10362 24552 10364
rect 24256 10310 24282 10362
rect 24282 10310 24312 10362
rect 24336 10310 24346 10362
rect 24346 10310 24392 10362
rect 24416 10310 24462 10362
rect 24462 10310 24472 10362
rect 24496 10310 24526 10362
rect 24526 10310 24552 10362
rect 24256 10308 24312 10310
rect 24336 10308 24392 10310
rect 24416 10308 24472 10310
rect 24496 10308 24552 10310
rect 27256 10362 27312 10364
rect 27336 10362 27392 10364
rect 27416 10362 27472 10364
rect 27496 10362 27552 10364
rect 27256 10310 27282 10362
rect 27282 10310 27312 10362
rect 27336 10310 27346 10362
rect 27346 10310 27392 10362
rect 27416 10310 27462 10362
rect 27462 10310 27472 10362
rect 27496 10310 27526 10362
rect 27526 10310 27552 10362
rect 27256 10308 27312 10310
rect 27336 10308 27392 10310
rect 27416 10308 27472 10310
rect 27496 10308 27552 10310
rect 22756 9818 22812 9820
rect 22836 9818 22892 9820
rect 22916 9818 22972 9820
rect 22996 9818 23052 9820
rect 22756 9766 22782 9818
rect 22782 9766 22812 9818
rect 22836 9766 22846 9818
rect 22846 9766 22892 9818
rect 22916 9766 22962 9818
rect 22962 9766 22972 9818
rect 22996 9766 23026 9818
rect 23026 9766 23052 9818
rect 22756 9764 22812 9766
rect 22836 9764 22892 9766
rect 22916 9764 22972 9766
rect 22996 9764 23052 9766
rect 25756 9818 25812 9820
rect 25836 9818 25892 9820
rect 25916 9818 25972 9820
rect 25996 9818 26052 9820
rect 25756 9766 25782 9818
rect 25782 9766 25812 9818
rect 25836 9766 25846 9818
rect 25846 9766 25892 9818
rect 25916 9766 25962 9818
rect 25962 9766 25972 9818
rect 25996 9766 26026 9818
rect 26026 9766 26052 9818
rect 25756 9764 25812 9766
rect 25836 9764 25892 9766
rect 25916 9764 25972 9766
rect 25996 9764 26052 9766
rect 24256 9274 24312 9276
rect 24336 9274 24392 9276
rect 24416 9274 24472 9276
rect 24496 9274 24552 9276
rect 24256 9222 24282 9274
rect 24282 9222 24312 9274
rect 24336 9222 24346 9274
rect 24346 9222 24392 9274
rect 24416 9222 24462 9274
rect 24462 9222 24472 9274
rect 24496 9222 24526 9274
rect 24526 9222 24552 9274
rect 24256 9220 24312 9222
rect 24336 9220 24392 9222
rect 24416 9220 24472 9222
rect 24496 9220 24552 9222
rect 27256 9274 27312 9276
rect 27336 9274 27392 9276
rect 27416 9274 27472 9276
rect 27496 9274 27552 9276
rect 27256 9222 27282 9274
rect 27282 9222 27312 9274
rect 27336 9222 27346 9274
rect 27346 9222 27392 9274
rect 27416 9222 27462 9274
rect 27462 9222 27472 9274
rect 27496 9222 27526 9274
rect 27526 9222 27552 9274
rect 27256 9220 27312 9222
rect 27336 9220 27392 9222
rect 27416 9220 27472 9222
rect 27496 9220 27552 9222
rect 22756 8730 22812 8732
rect 22836 8730 22892 8732
rect 22916 8730 22972 8732
rect 22996 8730 23052 8732
rect 22756 8678 22782 8730
rect 22782 8678 22812 8730
rect 22836 8678 22846 8730
rect 22846 8678 22892 8730
rect 22916 8678 22962 8730
rect 22962 8678 22972 8730
rect 22996 8678 23026 8730
rect 23026 8678 23052 8730
rect 22756 8676 22812 8678
rect 22836 8676 22892 8678
rect 22916 8676 22972 8678
rect 22996 8676 23052 8678
rect 25756 8730 25812 8732
rect 25836 8730 25892 8732
rect 25916 8730 25972 8732
rect 25996 8730 26052 8732
rect 25756 8678 25782 8730
rect 25782 8678 25812 8730
rect 25836 8678 25846 8730
rect 25846 8678 25892 8730
rect 25916 8678 25962 8730
rect 25962 8678 25972 8730
rect 25996 8678 26026 8730
rect 26026 8678 26052 8730
rect 25756 8676 25812 8678
rect 25836 8676 25892 8678
rect 25916 8676 25972 8678
rect 25996 8676 26052 8678
rect 24256 8186 24312 8188
rect 24336 8186 24392 8188
rect 24416 8186 24472 8188
rect 24496 8186 24552 8188
rect 24256 8134 24282 8186
rect 24282 8134 24312 8186
rect 24336 8134 24346 8186
rect 24346 8134 24392 8186
rect 24416 8134 24462 8186
rect 24462 8134 24472 8186
rect 24496 8134 24526 8186
rect 24526 8134 24552 8186
rect 24256 8132 24312 8134
rect 24336 8132 24392 8134
rect 24416 8132 24472 8134
rect 24496 8132 24552 8134
rect 27256 8186 27312 8188
rect 27336 8186 27392 8188
rect 27416 8186 27472 8188
rect 27496 8186 27552 8188
rect 27256 8134 27282 8186
rect 27282 8134 27312 8186
rect 27336 8134 27346 8186
rect 27346 8134 27392 8186
rect 27416 8134 27462 8186
rect 27462 8134 27472 8186
rect 27496 8134 27526 8186
rect 27526 8134 27552 8186
rect 27256 8132 27312 8134
rect 27336 8132 27392 8134
rect 27416 8132 27472 8134
rect 27496 8132 27552 8134
rect 22756 7642 22812 7644
rect 22836 7642 22892 7644
rect 22916 7642 22972 7644
rect 22996 7642 23052 7644
rect 22756 7590 22782 7642
rect 22782 7590 22812 7642
rect 22836 7590 22846 7642
rect 22846 7590 22892 7642
rect 22916 7590 22962 7642
rect 22962 7590 22972 7642
rect 22996 7590 23026 7642
rect 23026 7590 23052 7642
rect 22756 7588 22812 7590
rect 22836 7588 22892 7590
rect 22916 7588 22972 7590
rect 22996 7588 23052 7590
rect 25756 7642 25812 7644
rect 25836 7642 25892 7644
rect 25916 7642 25972 7644
rect 25996 7642 26052 7644
rect 25756 7590 25782 7642
rect 25782 7590 25812 7642
rect 25836 7590 25846 7642
rect 25846 7590 25892 7642
rect 25916 7590 25962 7642
rect 25962 7590 25972 7642
rect 25996 7590 26026 7642
rect 26026 7590 26052 7642
rect 25756 7588 25812 7590
rect 25836 7588 25892 7590
rect 25916 7588 25972 7590
rect 25996 7588 26052 7590
rect 24256 7098 24312 7100
rect 24336 7098 24392 7100
rect 24416 7098 24472 7100
rect 24496 7098 24552 7100
rect 24256 7046 24282 7098
rect 24282 7046 24312 7098
rect 24336 7046 24346 7098
rect 24346 7046 24392 7098
rect 24416 7046 24462 7098
rect 24462 7046 24472 7098
rect 24496 7046 24526 7098
rect 24526 7046 24552 7098
rect 24256 7044 24312 7046
rect 24336 7044 24392 7046
rect 24416 7044 24472 7046
rect 24496 7044 24552 7046
rect 27256 7098 27312 7100
rect 27336 7098 27392 7100
rect 27416 7098 27472 7100
rect 27496 7098 27552 7100
rect 27256 7046 27282 7098
rect 27282 7046 27312 7098
rect 27336 7046 27346 7098
rect 27346 7046 27392 7098
rect 27416 7046 27462 7098
rect 27462 7046 27472 7098
rect 27496 7046 27526 7098
rect 27526 7046 27552 7098
rect 27256 7044 27312 7046
rect 27336 7044 27392 7046
rect 27416 7044 27472 7046
rect 27496 7044 27552 7046
rect 21256 6010 21312 6012
rect 21336 6010 21392 6012
rect 21416 6010 21472 6012
rect 21496 6010 21552 6012
rect 21256 5958 21282 6010
rect 21282 5958 21312 6010
rect 21336 5958 21346 6010
rect 21346 5958 21392 6010
rect 21416 5958 21462 6010
rect 21462 5958 21472 6010
rect 21496 5958 21526 6010
rect 21526 5958 21552 6010
rect 21256 5956 21312 5958
rect 21336 5956 21392 5958
rect 21416 5956 21472 5958
rect 21496 5956 21552 5958
rect 22756 6554 22812 6556
rect 22836 6554 22892 6556
rect 22916 6554 22972 6556
rect 22996 6554 23052 6556
rect 22756 6502 22782 6554
rect 22782 6502 22812 6554
rect 22836 6502 22846 6554
rect 22846 6502 22892 6554
rect 22916 6502 22962 6554
rect 22962 6502 22972 6554
rect 22996 6502 23026 6554
rect 23026 6502 23052 6554
rect 22756 6500 22812 6502
rect 22836 6500 22892 6502
rect 22916 6500 22972 6502
rect 22996 6500 23052 6502
rect 25756 6554 25812 6556
rect 25836 6554 25892 6556
rect 25916 6554 25972 6556
rect 25996 6554 26052 6556
rect 25756 6502 25782 6554
rect 25782 6502 25812 6554
rect 25836 6502 25846 6554
rect 25846 6502 25892 6554
rect 25916 6502 25962 6554
rect 25962 6502 25972 6554
rect 25996 6502 26026 6554
rect 26026 6502 26052 6554
rect 25756 6500 25812 6502
rect 25836 6500 25892 6502
rect 25916 6500 25972 6502
rect 25996 6500 26052 6502
rect 24256 6010 24312 6012
rect 24336 6010 24392 6012
rect 24416 6010 24472 6012
rect 24496 6010 24552 6012
rect 24256 5958 24282 6010
rect 24282 5958 24312 6010
rect 24336 5958 24346 6010
rect 24346 5958 24392 6010
rect 24416 5958 24462 6010
rect 24462 5958 24472 6010
rect 24496 5958 24526 6010
rect 24526 5958 24552 6010
rect 24256 5956 24312 5958
rect 24336 5956 24392 5958
rect 24416 5956 24472 5958
rect 24496 5956 24552 5958
rect 27256 6010 27312 6012
rect 27336 6010 27392 6012
rect 27416 6010 27472 6012
rect 27496 6010 27552 6012
rect 27256 5958 27282 6010
rect 27282 5958 27312 6010
rect 27336 5958 27346 6010
rect 27346 5958 27392 6010
rect 27416 5958 27462 6010
rect 27462 5958 27472 6010
rect 27496 5958 27526 6010
rect 27526 5958 27552 6010
rect 27256 5956 27312 5958
rect 27336 5956 27392 5958
rect 27416 5956 27472 5958
rect 27496 5956 27552 5958
rect 22756 5466 22812 5468
rect 22836 5466 22892 5468
rect 22916 5466 22972 5468
rect 22996 5466 23052 5468
rect 22756 5414 22782 5466
rect 22782 5414 22812 5466
rect 22836 5414 22846 5466
rect 22846 5414 22892 5466
rect 22916 5414 22962 5466
rect 22962 5414 22972 5466
rect 22996 5414 23026 5466
rect 23026 5414 23052 5466
rect 22756 5412 22812 5414
rect 22836 5412 22892 5414
rect 22916 5412 22972 5414
rect 22996 5412 23052 5414
rect 25756 5466 25812 5468
rect 25836 5466 25892 5468
rect 25916 5466 25972 5468
rect 25996 5466 26052 5468
rect 25756 5414 25782 5466
rect 25782 5414 25812 5466
rect 25836 5414 25846 5466
rect 25846 5414 25892 5466
rect 25916 5414 25962 5466
rect 25962 5414 25972 5466
rect 25996 5414 26026 5466
rect 26026 5414 26052 5466
rect 25756 5412 25812 5414
rect 25836 5412 25892 5414
rect 25916 5412 25972 5414
rect 25996 5412 26052 5414
rect 19756 4378 19812 4380
rect 19836 4378 19892 4380
rect 19916 4378 19972 4380
rect 19996 4378 20052 4380
rect 19756 4326 19782 4378
rect 19782 4326 19812 4378
rect 19836 4326 19846 4378
rect 19846 4326 19892 4378
rect 19916 4326 19962 4378
rect 19962 4326 19972 4378
rect 19996 4326 20026 4378
rect 20026 4326 20052 4378
rect 19756 4324 19812 4326
rect 19836 4324 19892 4326
rect 19916 4324 19972 4326
rect 19996 4324 20052 4326
rect 21256 4922 21312 4924
rect 21336 4922 21392 4924
rect 21416 4922 21472 4924
rect 21496 4922 21552 4924
rect 21256 4870 21282 4922
rect 21282 4870 21312 4922
rect 21336 4870 21346 4922
rect 21346 4870 21392 4922
rect 21416 4870 21462 4922
rect 21462 4870 21472 4922
rect 21496 4870 21526 4922
rect 21526 4870 21552 4922
rect 21256 4868 21312 4870
rect 21336 4868 21392 4870
rect 21416 4868 21472 4870
rect 21496 4868 21552 4870
rect 24256 4922 24312 4924
rect 24336 4922 24392 4924
rect 24416 4922 24472 4924
rect 24496 4922 24552 4924
rect 24256 4870 24282 4922
rect 24282 4870 24312 4922
rect 24336 4870 24346 4922
rect 24346 4870 24392 4922
rect 24416 4870 24462 4922
rect 24462 4870 24472 4922
rect 24496 4870 24526 4922
rect 24526 4870 24552 4922
rect 24256 4868 24312 4870
rect 24336 4868 24392 4870
rect 24416 4868 24472 4870
rect 24496 4868 24552 4870
rect 27256 4922 27312 4924
rect 27336 4922 27392 4924
rect 27416 4922 27472 4924
rect 27496 4922 27552 4924
rect 27256 4870 27282 4922
rect 27282 4870 27312 4922
rect 27336 4870 27346 4922
rect 27346 4870 27392 4922
rect 27416 4870 27462 4922
rect 27462 4870 27472 4922
rect 27496 4870 27526 4922
rect 27526 4870 27552 4922
rect 27256 4868 27312 4870
rect 27336 4868 27392 4870
rect 27416 4868 27472 4870
rect 27496 4868 27552 4870
rect 22756 4378 22812 4380
rect 22836 4378 22892 4380
rect 22916 4378 22972 4380
rect 22996 4378 23052 4380
rect 22756 4326 22782 4378
rect 22782 4326 22812 4378
rect 22836 4326 22846 4378
rect 22846 4326 22892 4378
rect 22916 4326 22962 4378
rect 22962 4326 22972 4378
rect 22996 4326 23026 4378
rect 23026 4326 23052 4378
rect 22756 4324 22812 4326
rect 22836 4324 22892 4326
rect 22916 4324 22972 4326
rect 22996 4324 23052 4326
rect 25756 4378 25812 4380
rect 25836 4378 25892 4380
rect 25916 4378 25972 4380
rect 25996 4378 26052 4380
rect 25756 4326 25782 4378
rect 25782 4326 25812 4378
rect 25836 4326 25846 4378
rect 25846 4326 25892 4378
rect 25916 4326 25962 4378
rect 25962 4326 25972 4378
rect 25996 4326 26026 4378
rect 26026 4326 26052 4378
rect 25756 4324 25812 4326
rect 25836 4324 25892 4326
rect 25916 4324 25972 4326
rect 25996 4324 26052 4326
rect 18256 3834 18312 3836
rect 18336 3834 18392 3836
rect 18416 3834 18472 3836
rect 18496 3834 18552 3836
rect 18256 3782 18282 3834
rect 18282 3782 18312 3834
rect 18336 3782 18346 3834
rect 18346 3782 18392 3834
rect 18416 3782 18462 3834
rect 18462 3782 18472 3834
rect 18496 3782 18526 3834
rect 18526 3782 18552 3834
rect 18256 3780 18312 3782
rect 18336 3780 18392 3782
rect 18416 3780 18472 3782
rect 18496 3780 18552 3782
rect 16756 3290 16812 3292
rect 16836 3290 16892 3292
rect 16916 3290 16972 3292
rect 16996 3290 17052 3292
rect 16756 3238 16782 3290
rect 16782 3238 16812 3290
rect 16836 3238 16846 3290
rect 16846 3238 16892 3290
rect 16916 3238 16962 3290
rect 16962 3238 16972 3290
rect 16996 3238 17026 3290
rect 17026 3238 17052 3290
rect 16756 3236 16812 3238
rect 16836 3236 16892 3238
rect 16916 3236 16972 3238
rect 16996 3236 17052 3238
rect 15256 2746 15312 2748
rect 15336 2746 15392 2748
rect 15416 2746 15472 2748
rect 15496 2746 15552 2748
rect 15256 2694 15282 2746
rect 15282 2694 15312 2746
rect 15336 2694 15346 2746
rect 15346 2694 15392 2746
rect 15416 2694 15462 2746
rect 15462 2694 15472 2746
rect 15496 2694 15526 2746
rect 15526 2694 15552 2746
rect 15256 2692 15312 2694
rect 15336 2692 15392 2694
rect 15416 2692 15472 2694
rect 15496 2692 15552 2694
rect 18256 2746 18312 2748
rect 18336 2746 18392 2748
rect 18416 2746 18472 2748
rect 18496 2746 18552 2748
rect 18256 2694 18282 2746
rect 18282 2694 18312 2746
rect 18336 2694 18346 2746
rect 18346 2694 18392 2746
rect 18416 2694 18462 2746
rect 18462 2694 18472 2746
rect 18496 2694 18526 2746
rect 18526 2694 18552 2746
rect 18256 2692 18312 2694
rect 18336 2692 18392 2694
rect 18416 2692 18472 2694
rect 18496 2692 18552 2694
rect 21256 3834 21312 3836
rect 21336 3834 21392 3836
rect 21416 3834 21472 3836
rect 21496 3834 21552 3836
rect 21256 3782 21282 3834
rect 21282 3782 21312 3834
rect 21336 3782 21346 3834
rect 21346 3782 21392 3834
rect 21416 3782 21462 3834
rect 21462 3782 21472 3834
rect 21496 3782 21526 3834
rect 21526 3782 21552 3834
rect 21256 3780 21312 3782
rect 21336 3780 21392 3782
rect 21416 3780 21472 3782
rect 21496 3780 21552 3782
rect 24256 3834 24312 3836
rect 24336 3834 24392 3836
rect 24416 3834 24472 3836
rect 24496 3834 24552 3836
rect 24256 3782 24282 3834
rect 24282 3782 24312 3834
rect 24336 3782 24346 3834
rect 24346 3782 24392 3834
rect 24416 3782 24462 3834
rect 24462 3782 24472 3834
rect 24496 3782 24526 3834
rect 24526 3782 24552 3834
rect 24256 3780 24312 3782
rect 24336 3780 24392 3782
rect 24416 3780 24472 3782
rect 24496 3780 24552 3782
rect 27256 3834 27312 3836
rect 27336 3834 27392 3836
rect 27416 3834 27472 3836
rect 27496 3834 27552 3836
rect 27256 3782 27282 3834
rect 27282 3782 27312 3834
rect 27336 3782 27346 3834
rect 27346 3782 27392 3834
rect 27416 3782 27462 3834
rect 27462 3782 27472 3834
rect 27496 3782 27526 3834
rect 27526 3782 27552 3834
rect 27256 3780 27312 3782
rect 27336 3780 27392 3782
rect 27416 3780 27472 3782
rect 27496 3780 27552 3782
rect 19756 3290 19812 3292
rect 19836 3290 19892 3292
rect 19916 3290 19972 3292
rect 19996 3290 20052 3292
rect 19756 3238 19782 3290
rect 19782 3238 19812 3290
rect 19836 3238 19846 3290
rect 19846 3238 19892 3290
rect 19916 3238 19962 3290
rect 19962 3238 19972 3290
rect 19996 3238 20026 3290
rect 20026 3238 20052 3290
rect 19756 3236 19812 3238
rect 19836 3236 19892 3238
rect 19916 3236 19972 3238
rect 19996 3236 20052 3238
rect 22756 3290 22812 3292
rect 22836 3290 22892 3292
rect 22916 3290 22972 3292
rect 22996 3290 23052 3292
rect 22756 3238 22782 3290
rect 22782 3238 22812 3290
rect 22836 3238 22846 3290
rect 22846 3238 22892 3290
rect 22916 3238 22962 3290
rect 22962 3238 22972 3290
rect 22996 3238 23026 3290
rect 23026 3238 23052 3290
rect 22756 3236 22812 3238
rect 22836 3236 22892 3238
rect 22916 3236 22972 3238
rect 22996 3236 23052 3238
rect 25756 3290 25812 3292
rect 25836 3290 25892 3292
rect 25916 3290 25972 3292
rect 25996 3290 26052 3292
rect 25756 3238 25782 3290
rect 25782 3238 25812 3290
rect 25836 3238 25846 3290
rect 25846 3238 25892 3290
rect 25916 3238 25962 3290
rect 25962 3238 25972 3290
rect 25996 3238 26026 3290
rect 26026 3238 26052 3290
rect 25756 3236 25812 3238
rect 25836 3236 25892 3238
rect 25916 3236 25972 3238
rect 25996 3236 26052 3238
rect 21256 2746 21312 2748
rect 21336 2746 21392 2748
rect 21416 2746 21472 2748
rect 21496 2746 21552 2748
rect 21256 2694 21282 2746
rect 21282 2694 21312 2746
rect 21336 2694 21346 2746
rect 21346 2694 21392 2746
rect 21416 2694 21462 2746
rect 21462 2694 21472 2746
rect 21496 2694 21526 2746
rect 21526 2694 21552 2746
rect 21256 2692 21312 2694
rect 21336 2692 21392 2694
rect 21416 2692 21472 2694
rect 21496 2692 21552 2694
rect 24256 2746 24312 2748
rect 24336 2746 24392 2748
rect 24416 2746 24472 2748
rect 24496 2746 24552 2748
rect 24256 2694 24282 2746
rect 24282 2694 24312 2746
rect 24336 2694 24346 2746
rect 24346 2694 24392 2746
rect 24416 2694 24462 2746
rect 24462 2694 24472 2746
rect 24496 2694 24526 2746
rect 24526 2694 24552 2746
rect 24256 2692 24312 2694
rect 24336 2692 24392 2694
rect 24416 2692 24472 2694
rect 24496 2692 24552 2694
rect 27256 2746 27312 2748
rect 27336 2746 27392 2748
rect 27416 2746 27472 2748
rect 27496 2746 27552 2748
rect 27256 2694 27282 2746
rect 27282 2694 27312 2746
rect 27336 2694 27346 2746
rect 27346 2694 27392 2746
rect 27416 2694 27462 2746
rect 27462 2694 27472 2746
rect 27496 2694 27526 2746
rect 27526 2694 27552 2746
rect 27256 2692 27312 2694
rect 27336 2692 27392 2694
rect 27416 2692 27472 2694
rect 27496 2692 27552 2694
rect 10756 2202 10812 2204
rect 10836 2202 10892 2204
rect 10916 2202 10972 2204
rect 10996 2202 11052 2204
rect 10756 2150 10782 2202
rect 10782 2150 10812 2202
rect 10836 2150 10846 2202
rect 10846 2150 10892 2202
rect 10916 2150 10962 2202
rect 10962 2150 10972 2202
rect 10996 2150 11026 2202
rect 11026 2150 11052 2202
rect 10756 2148 10812 2150
rect 10836 2148 10892 2150
rect 10916 2148 10972 2150
rect 10996 2148 11052 2150
rect 13756 2202 13812 2204
rect 13836 2202 13892 2204
rect 13916 2202 13972 2204
rect 13996 2202 14052 2204
rect 13756 2150 13782 2202
rect 13782 2150 13812 2202
rect 13836 2150 13846 2202
rect 13846 2150 13892 2202
rect 13916 2150 13962 2202
rect 13962 2150 13972 2202
rect 13996 2150 14026 2202
rect 14026 2150 14052 2202
rect 13756 2148 13812 2150
rect 13836 2148 13892 2150
rect 13916 2148 13972 2150
rect 13996 2148 14052 2150
rect 16756 2202 16812 2204
rect 16836 2202 16892 2204
rect 16916 2202 16972 2204
rect 16996 2202 17052 2204
rect 16756 2150 16782 2202
rect 16782 2150 16812 2202
rect 16836 2150 16846 2202
rect 16846 2150 16892 2202
rect 16916 2150 16962 2202
rect 16962 2150 16972 2202
rect 16996 2150 17026 2202
rect 17026 2150 17052 2202
rect 16756 2148 16812 2150
rect 16836 2148 16892 2150
rect 16916 2148 16972 2150
rect 16996 2148 17052 2150
rect 19756 2202 19812 2204
rect 19836 2202 19892 2204
rect 19916 2202 19972 2204
rect 19996 2202 20052 2204
rect 19756 2150 19782 2202
rect 19782 2150 19812 2202
rect 19836 2150 19846 2202
rect 19846 2150 19892 2202
rect 19916 2150 19962 2202
rect 19962 2150 19972 2202
rect 19996 2150 20026 2202
rect 20026 2150 20052 2202
rect 19756 2148 19812 2150
rect 19836 2148 19892 2150
rect 19916 2148 19972 2150
rect 19996 2148 20052 2150
rect 22756 2202 22812 2204
rect 22836 2202 22892 2204
rect 22916 2202 22972 2204
rect 22996 2202 23052 2204
rect 22756 2150 22782 2202
rect 22782 2150 22812 2202
rect 22836 2150 22846 2202
rect 22846 2150 22892 2202
rect 22916 2150 22962 2202
rect 22962 2150 22972 2202
rect 22996 2150 23026 2202
rect 23026 2150 23052 2202
rect 22756 2148 22812 2150
rect 22836 2148 22892 2150
rect 22916 2148 22972 2150
rect 22996 2148 23052 2150
rect 25756 2202 25812 2204
rect 25836 2202 25892 2204
rect 25916 2202 25972 2204
rect 25996 2202 26052 2204
rect 25756 2150 25782 2202
rect 25782 2150 25812 2202
rect 25836 2150 25846 2202
rect 25846 2150 25892 2202
rect 25916 2150 25962 2202
rect 25962 2150 25972 2202
rect 25996 2150 26026 2202
rect 26026 2150 26052 2202
rect 25756 2148 25812 2150
rect 25836 2148 25892 2150
rect 25916 2148 25972 2150
rect 25996 2148 26052 2150
<< metal3 >>
rect 1744 29408 2064 29409
rect 1744 29344 1752 29408
rect 1816 29344 1832 29408
rect 1896 29344 1912 29408
rect 1976 29344 1992 29408
rect 2056 29344 2064 29408
rect 1744 29343 2064 29344
rect 4744 29408 5064 29409
rect 4744 29344 4752 29408
rect 4816 29344 4832 29408
rect 4896 29344 4912 29408
rect 4976 29344 4992 29408
rect 5056 29344 5064 29408
rect 4744 29343 5064 29344
rect 7744 29408 8064 29409
rect 7744 29344 7752 29408
rect 7816 29344 7832 29408
rect 7896 29344 7912 29408
rect 7976 29344 7992 29408
rect 8056 29344 8064 29408
rect 7744 29343 8064 29344
rect 10744 29408 11064 29409
rect 10744 29344 10752 29408
rect 10816 29344 10832 29408
rect 10896 29344 10912 29408
rect 10976 29344 10992 29408
rect 11056 29344 11064 29408
rect 10744 29343 11064 29344
rect 13744 29408 14064 29409
rect 13744 29344 13752 29408
rect 13816 29344 13832 29408
rect 13896 29344 13912 29408
rect 13976 29344 13992 29408
rect 14056 29344 14064 29408
rect 13744 29343 14064 29344
rect 16744 29408 17064 29409
rect 16744 29344 16752 29408
rect 16816 29344 16832 29408
rect 16896 29344 16912 29408
rect 16976 29344 16992 29408
rect 17056 29344 17064 29408
rect 16744 29343 17064 29344
rect 19744 29408 20064 29409
rect 19744 29344 19752 29408
rect 19816 29344 19832 29408
rect 19896 29344 19912 29408
rect 19976 29344 19992 29408
rect 20056 29344 20064 29408
rect 19744 29343 20064 29344
rect 22744 29408 23064 29409
rect 22744 29344 22752 29408
rect 22816 29344 22832 29408
rect 22896 29344 22912 29408
rect 22976 29344 22992 29408
rect 23056 29344 23064 29408
rect 22744 29343 23064 29344
rect 25744 29408 26064 29409
rect 25744 29344 25752 29408
rect 25816 29344 25832 29408
rect 25896 29344 25912 29408
rect 25976 29344 25992 29408
rect 26056 29344 26064 29408
rect 25744 29343 26064 29344
rect 3244 28864 3564 28865
rect 3244 28800 3252 28864
rect 3316 28800 3332 28864
rect 3396 28800 3412 28864
rect 3476 28800 3492 28864
rect 3556 28800 3564 28864
rect 3244 28799 3564 28800
rect 6244 28864 6564 28865
rect 6244 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6412 28864
rect 6476 28800 6492 28864
rect 6556 28800 6564 28864
rect 6244 28799 6564 28800
rect 9244 28864 9564 28865
rect 9244 28800 9252 28864
rect 9316 28800 9332 28864
rect 9396 28800 9412 28864
rect 9476 28800 9492 28864
rect 9556 28800 9564 28864
rect 9244 28799 9564 28800
rect 12244 28864 12564 28865
rect 12244 28800 12252 28864
rect 12316 28800 12332 28864
rect 12396 28800 12412 28864
rect 12476 28800 12492 28864
rect 12556 28800 12564 28864
rect 12244 28799 12564 28800
rect 15244 28864 15564 28865
rect 15244 28800 15252 28864
rect 15316 28800 15332 28864
rect 15396 28800 15412 28864
rect 15476 28800 15492 28864
rect 15556 28800 15564 28864
rect 15244 28799 15564 28800
rect 18244 28864 18564 28865
rect 18244 28800 18252 28864
rect 18316 28800 18332 28864
rect 18396 28800 18412 28864
rect 18476 28800 18492 28864
rect 18556 28800 18564 28864
rect 18244 28799 18564 28800
rect 21244 28864 21564 28865
rect 21244 28800 21252 28864
rect 21316 28800 21332 28864
rect 21396 28800 21412 28864
rect 21476 28800 21492 28864
rect 21556 28800 21564 28864
rect 21244 28799 21564 28800
rect 24244 28864 24564 28865
rect 24244 28800 24252 28864
rect 24316 28800 24332 28864
rect 24396 28800 24412 28864
rect 24476 28800 24492 28864
rect 24556 28800 24564 28864
rect 24244 28799 24564 28800
rect 27244 28864 27564 28865
rect 27244 28800 27252 28864
rect 27316 28800 27332 28864
rect 27396 28800 27412 28864
rect 27476 28800 27492 28864
rect 27556 28800 27564 28864
rect 27244 28799 27564 28800
rect 1744 28320 2064 28321
rect 1744 28256 1752 28320
rect 1816 28256 1832 28320
rect 1896 28256 1912 28320
rect 1976 28256 1992 28320
rect 2056 28256 2064 28320
rect 1744 28255 2064 28256
rect 4744 28320 5064 28321
rect 4744 28256 4752 28320
rect 4816 28256 4832 28320
rect 4896 28256 4912 28320
rect 4976 28256 4992 28320
rect 5056 28256 5064 28320
rect 4744 28255 5064 28256
rect 7744 28320 8064 28321
rect 7744 28256 7752 28320
rect 7816 28256 7832 28320
rect 7896 28256 7912 28320
rect 7976 28256 7992 28320
rect 8056 28256 8064 28320
rect 7744 28255 8064 28256
rect 10744 28320 11064 28321
rect 10744 28256 10752 28320
rect 10816 28256 10832 28320
rect 10896 28256 10912 28320
rect 10976 28256 10992 28320
rect 11056 28256 11064 28320
rect 10744 28255 11064 28256
rect 13744 28320 14064 28321
rect 13744 28256 13752 28320
rect 13816 28256 13832 28320
rect 13896 28256 13912 28320
rect 13976 28256 13992 28320
rect 14056 28256 14064 28320
rect 13744 28255 14064 28256
rect 16744 28320 17064 28321
rect 16744 28256 16752 28320
rect 16816 28256 16832 28320
rect 16896 28256 16912 28320
rect 16976 28256 16992 28320
rect 17056 28256 17064 28320
rect 16744 28255 17064 28256
rect 19744 28320 20064 28321
rect 19744 28256 19752 28320
rect 19816 28256 19832 28320
rect 19896 28256 19912 28320
rect 19976 28256 19992 28320
rect 20056 28256 20064 28320
rect 19744 28255 20064 28256
rect 22744 28320 23064 28321
rect 22744 28256 22752 28320
rect 22816 28256 22832 28320
rect 22896 28256 22912 28320
rect 22976 28256 22992 28320
rect 23056 28256 23064 28320
rect 22744 28255 23064 28256
rect 25744 28320 26064 28321
rect 25744 28256 25752 28320
rect 25816 28256 25832 28320
rect 25896 28256 25912 28320
rect 25976 28256 25992 28320
rect 26056 28256 26064 28320
rect 25744 28255 26064 28256
rect 3244 27776 3564 27777
rect 3244 27712 3252 27776
rect 3316 27712 3332 27776
rect 3396 27712 3412 27776
rect 3476 27712 3492 27776
rect 3556 27712 3564 27776
rect 3244 27711 3564 27712
rect 6244 27776 6564 27777
rect 6244 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6412 27776
rect 6476 27712 6492 27776
rect 6556 27712 6564 27776
rect 6244 27711 6564 27712
rect 9244 27776 9564 27777
rect 9244 27712 9252 27776
rect 9316 27712 9332 27776
rect 9396 27712 9412 27776
rect 9476 27712 9492 27776
rect 9556 27712 9564 27776
rect 9244 27711 9564 27712
rect 12244 27776 12564 27777
rect 12244 27712 12252 27776
rect 12316 27712 12332 27776
rect 12396 27712 12412 27776
rect 12476 27712 12492 27776
rect 12556 27712 12564 27776
rect 12244 27711 12564 27712
rect 15244 27776 15564 27777
rect 15244 27712 15252 27776
rect 15316 27712 15332 27776
rect 15396 27712 15412 27776
rect 15476 27712 15492 27776
rect 15556 27712 15564 27776
rect 15244 27711 15564 27712
rect 18244 27776 18564 27777
rect 18244 27712 18252 27776
rect 18316 27712 18332 27776
rect 18396 27712 18412 27776
rect 18476 27712 18492 27776
rect 18556 27712 18564 27776
rect 18244 27711 18564 27712
rect 21244 27776 21564 27777
rect 21244 27712 21252 27776
rect 21316 27712 21332 27776
rect 21396 27712 21412 27776
rect 21476 27712 21492 27776
rect 21556 27712 21564 27776
rect 21244 27711 21564 27712
rect 24244 27776 24564 27777
rect 24244 27712 24252 27776
rect 24316 27712 24332 27776
rect 24396 27712 24412 27776
rect 24476 27712 24492 27776
rect 24556 27712 24564 27776
rect 24244 27711 24564 27712
rect 27244 27776 27564 27777
rect 27244 27712 27252 27776
rect 27316 27712 27332 27776
rect 27396 27712 27412 27776
rect 27476 27712 27492 27776
rect 27556 27712 27564 27776
rect 27244 27711 27564 27712
rect 0 27344 800 27464
rect 1744 27232 2064 27233
rect 1744 27168 1752 27232
rect 1816 27168 1832 27232
rect 1896 27168 1912 27232
rect 1976 27168 1992 27232
rect 2056 27168 2064 27232
rect 1744 27167 2064 27168
rect 4744 27232 5064 27233
rect 4744 27168 4752 27232
rect 4816 27168 4832 27232
rect 4896 27168 4912 27232
rect 4976 27168 4992 27232
rect 5056 27168 5064 27232
rect 4744 27167 5064 27168
rect 7744 27232 8064 27233
rect 7744 27168 7752 27232
rect 7816 27168 7832 27232
rect 7896 27168 7912 27232
rect 7976 27168 7992 27232
rect 8056 27168 8064 27232
rect 7744 27167 8064 27168
rect 10744 27232 11064 27233
rect 10744 27168 10752 27232
rect 10816 27168 10832 27232
rect 10896 27168 10912 27232
rect 10976 27168 10992 27232
rect 11056 27168 11064 27232
rect 10744 27167 11064 27168
rect 13744 27232 14064 27233
rect 13744 27168 13752 27232
rect 13816 27168 13832 27232
rect 13896 27168 13912 27232
rect 13976 27168 13992 27232
rect 14056 27168 14064 27232
rect 13744 27167 14064 27168
rect 16744 27232 17064 27233
rect 16744 27168 16752 27232
rect 16816 27168 16832 27232
rect 16896 27168 16912 27232
rect 16976 27168 16992 27232
rect 17056 27168 17064 27232
rect 16744 27167 17064 27168
rect 19744 27232 20064 27233
rect 19744 27168 19752 27232
rect 19816 27168 19832 27232
rect 19896 27168 19912 27232
rect 19976 27168 19992 27232
rect 20056 27168 20064 27232
rect 19744 27167 20064 27168
rect 22744 27232 23064 27233
rect 22744 27168 22752 27232
rect 22816 27168 22832 27232
rect 22896 27168 22912 27232
rect 22976 27168 22992 27232
rect 23056 27168 23064 27232
rect 22744 27167 23064 27168
rect 25744 27232 26064 27233
rect 25744 27168 25752 27232
rect 25816 27168 25832 27232
rect 25896 27168 25912 27232
rect 25976 27168 25992 27232
rect 26056 27168 26064 27232
rect 25744 27167 26064 27168
rect 3244 26688 3564 26689
rect 3244 26624 3252 26688
rect 3316 26624 3332 26688
rect 3396 26624 3412 26688
rect 3476 26624 3492 26688
rect 3556 26624 3564 26688
rect 3244 26623 3564 26624
rect 6244 26688 6564 26689
rect 6244 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6412 26688
rect 6476 26624 6492 26688
rect 6556 26624 6564 26688
rect 6244 26623 6564 26624
rect 9244 26688 9564 26689
rect 9244 26624 9252 26688
rect 9316 26624 9332 26688
rect 9396 26624 9412 26688
rect 9476 26624 9492 26688
rect 9556 26624 9564 26688
rect 9244 26623 9564 26624
rect 12244 26688 12564 26689
rect 12244 26624 12252 26688
rect 12316 26624 12332 26688
rect 12396 26624 12412 26688
rect 12476 26624 12492 26688
rect 12556 26624 12564 26688
rect 12244 26623 12564 26624
rect 15244 26688 15564 26689
rect 15244 26624 15252 26688
rect 15316 26624 15332 26688
rect 15396 26624 15412 26688
rect 15476 26624 15492 26688
rect 15556 26624 15564 26688
rect 15244 26623 15564 26624
rect 18244 26688 18564 26689
rect 18244 26624 18252 26688
rect 18316 26624 18332 26688
rect 18396 26624 18412 26688
rect 18476 26624 18492 26688
rect 18556 26624 18564 26688
rect 18244 26623 18564 26624
rect 21244 26688 21564 26689
rect 21244 26624 21252 26688
rect 21316 26624 21332 26688
rect 21396 26624 21412 26688
rect 21476 26624 21492 26688
rect 21556 26624 21564 26688
rect 21244 26623 21564 26624
rect 24244 26688 24564 26689
rect 24244 26624 24252 26688
rect 24316 26624 24332 26688
rect 24396 26624 24412 26688
rect 24476 26624 24492 26688
rect 24556 26624 24564 26688
rect 24244 26623 24564 26624
rect 27244 26688 27564 26689
rect 27244 26624 27252 26688
rect 27316 26624 27332 26688
rect 27396 26624 27412 26688
rect 27476 26624 27492 26688
rect 27556 26624 27564 26688
rect 27244 26623 27564 26624
rect 1744 26144 2064 26145
rect 1744 26080 1752 26144
rect 1816 26080 1832 26144
rect 1896 26080 1912 26144
rect 1976 26080 1992 26144
rect 2056 26080 2064 26144
rect 1744 26079 2064 26080
rect 4744 26144 5064 26145
rect 4744 26080 4752 26144
rect 4816 26080 4832 26144
rect 4896 26080 4912 26144
rect 4976 26080 4992 26144
rect 5056 26080 5064 26144
rect 4744 26079 5064 26080
rect 7744 26144 8064 26145
rect 7744 26080 7752 26144
rect 7816 26080 7832 26144
rect 7896 26080 7912 26144
rect 7976 26080 7992 26144
rect 8056 26080 8064 26144
rect 7744 26079 8064 26080
rect 10744 26144 11064 26145
rect 10744 26080 10752 26144
rect 10816 26080 10832 26144
rect 10896 26080 10912 26144
rect 10976 26080 10992 26144
rect 11056 26080 11064 26144
rect 10744 26079 11064 26080
rect 13744 26144 14064 26145
rect 13744 26080 13752 26144
rect 13816 26080 13832 26144
rect 13896 26080 13912 26144
rect 13976 26080 13992 26144
rect 14056 26080 14064 26144
rect 13744 26079 14064 26080
rect 16744 26144 17064 26145
rect 16744 26080 16752 26144
rect 16816 26080 16832 26144
rect 16896 26080 16912 26144
rect 16976 26080 16992 26144
rect 17056 26080 17064 26144
rect 16744 26079 17064 26080
rect 19744 26144 20064 26145
rect 19744 26080 19752 26144
rect 19816 26080 19832 26144
rect 19896 26080 19912 26144
rect 19976 26080 19992 26144
rect 20056 26080 20064 26144
rect 19744 26079 20064 26080
rect 22744 26144 23064 26145
rect 22744 26080 22752 26144
rect 22816 26080 22832 26144
rect 22896 26080 22912 26144
rect 22976 26080 22992 26144
rect 23056 26080 23064 26144
rect 22744 26079 23064 26080
rect 25744 26144 26064 26145
rect 25744 26080 25752 26144
rect 25816 26080 25832 26144
rect 25896 26080 25912 26144
rect 25976 26080 25992 26144
rect 26056 26080 26064 26144
rect 25744 26079 26064 26080
rect 3244 25600 3564 25601
rect 3244 25536 3252 25600
rect 3316 25536 3332 25600
rect 3396 25536 3412 25600
rect 3476 25536 3492 25600
rect 3556 25536 3564 25600
rect 3244 25535 3564 25536
rect 6244 25600 6564 25601
rect 6244 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6412 25600
rect 6476 25536 6492 25600
rect 6556 25536 6564 25600
rect 6244 25535 6564 25536
rect 9244 25600 9564 25601
rect 9244 25536 9252 25600
rect 9316 25536 9332 25600
rect 9396 25536 9412 25600
rect 9476 25536 9492 25600
rect 9556 25536 9564 25600
rect 9244 25535 9564 25536
rect 12244 25600 12564 25601
rect 12244 25536 12252 25600
rect 12316 25536 12332 25600
rect 12396 25536 12412 25600
rect 12476 25536 12492 25600
rect 12556 25536 12564 25600
rect 12244 25535 12564 25536
rect 15244 25600 15564 25601
rect 15244 25536 15252 25600
rect 15316 25536 15332 25600
rect 15396 25536 15412 25600
rect 15476 25536 15492 25600
rect 15556 25536 15564 25600
rect 15244 25535 15564 25536
rect 18244 25600 18564 25601
rect 18244 25536 18252 25600
rect 18316 25536 18332 25600
rect 18396 25536 18412 25600
rect 18476 25536 18492 25600
rect 18556 25536 18564 25600
rect 18244 25535 18564 25536
rect 21244 25600 21564 25601
rect 21244 25536 21252 25600
rect 21316 25536 21332 25600
rect 21396 25536 21412 25600
rect 21476 25536 21492 25600
rect 21556 25536 21564 25600
rect 21244 25535 21564 25536
rect 24244 25600 24564 25601
rect 24244 25536 24252 25600
rect 24316 25536 24332 25600
rect 24396 25536 24412 25600
rect 24476 25536 24492 25600
rect 24556 25536 24564 25600
rect 24244 25535 24564 25536
rect 27244 25600 27564 25601
rect 27244 25536 27252 25600
rect 27316 25536 27332 25600
rect 27396 25536 27412 25600
rect 27476 25536 27492 25600
rect 27556 25536 27564 25600
rect 27244 25535 27564 25536
rect 1744 25056 2064 25057
rect 1744 24992 1752 25056
rect 1816 24992 1832 25056
rect 1896 24992 1912 25056
rect 1976 24992 1992 25056
rect 2056 24992 2064 25056
rect 1744 24991 2064 24992
rect 4744 25056 5064 25057
rect 4744 24992 4752 25056
rect 4816 24992 4832 25056
rect 4896 24992 4912 25056
rect 4976 24992 4992 25056
rect 5056 24992 5064 25056
rect 4744 24991 5064 24992
rect 7744 25056 8064 25057
rect 7744 24992 7752 25056
rect 7816 24992 7832 25056
rect 7896 24992 7912 25056
rect 7976 24992 7992 25056
rect 8056 24992 8064 25056
rect 7744 24991 8064 24992
rect 10744 25056 11064 25057
rect 10744 24992 10752 25056
rect 10816 24992 10832 25056
rect 10896 24992 10912 25056
rect 10976 24992 10992 25056
rect 11056 24992 11064 25056
rect 10744 24991 11064 24992
rect 13744 25056 14064 25057
rect 13744 24992 13752 25056
rect 13816 24992 13832 25056
rect 13896 24992 13912 25056
rect 13976 24992 13992 25056
rect 14056 24992 14064 25056
rect 13744 24991 14064 24992
rect 16744 25056 17064 25057
rect 16744 24992 16752 25056
rect 16816 24992 16832 25056
rect 16896 24992 16912 25056
rect 16976 24992 16992 25056
rect 17056 24992 17064 25056
rect 16744 24991 17064 24992
rect 19744 25056 20064 25057
rect 19744 24992 19752 25056
rect 19816 24992 19832 25056
rect 19896 24992 19912 25056
rect 19976 24992 19992 25056
rect 20056 24992 20064 25056
rect 19744 24991 20064 24992
rect 22744 25056 23064 25057
rect 22744 24992 22752 25056
rect 22816 24992 22832 25056
rect 22896 24992 22912 25056
rect 22976 24992 22992 25056
rect 23056 24992 23064 25056
rect 22744 24991 23064 24992
rect 25744 25056 26064 25057
rect 25744 24992 25752 25056
rect 25816 24992 25832 25056
rect 25896 24992 25912 25056
rect 25976 24992 25992 25056
rect 26056 24992 26064 25056
rect 25744 24991 26064 24992
rect 28727 24624 29527 24744
rect 3244 24512 3564 24513
rect 3244 24448 3252 24512
rect 3316 24448 3332 24512
rect 3396 24448 3412 24512
rect 3476 24448 3492 24512
rect 3556 24448 3564 24512
rect 3244 24447 3564 24448
rect 6244 24512 6564 24513
rect 6244 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6412 24512
rect 6476 24448 6492 24512
rect 6556 24448 6564 24512
rect 6244 24447 6564 24448
rect 9244 24512 9564 24513
rect 9244 24448 9252 24512
rect 9316 24448 9332 24512
rect 9396 24448 9412 24512
rect 9476 24448 9492 24512
rect 9556 24448 9564 24512
rect 9244 24447 9564 24448
rect 12244 24512 12564 24513
rect 12244 24448 12252 24512
rect 12316 24448 12332 24512
rect 12396 24448 12412 24512
rect 12476 24448 12492 24512
rect 12556 24448 12564 24512
rect 12244 24447 12564 24448
rect 15244 24512 15564 24513
rect 15244 24448 15252 24512
rect 15316 24448 15332 24512
rect 15396 24448 15412 24512
rect 15476 24448 15492 24512
rect 15556 24448 15564 24512
rect 15244 24447 15564 24448
rect 18244 24512 18564 24513
rect 18244 24448 18252 24512
rect 18316 24448 18332 24512
rect 18396 24448 18412 24512
rect 18476 24448 18492 24512
rect 18556 24448 18564 24512
rect 18244 24447 18564 24448
rect 21244 24512 21564 24513
rect 21244 24448 21252 24512
rect 21316 24448 21332 24512
rect 21396 24448 21412 24512
rect 21476 24448 21492 24512
rect 21556 24448 21564 24512
rect 21244 24447 21564 24448
rect 24244 24512 24564 24513
rect 24244 24448 24252 24512
rect 24316 24448 24332 24512
rect 24396 24448 24412 24512
rect 24476 24448 24492 24512
rect 24556 24448 24564 24512
rect 24244 24447 24564 24448
rect 27244 24512 27564 24513
rect 27244 24448 27252 24512
rect 27316 24448 27332 24512
rect 27396 24448 27412 24512
rect 27476 24448 27492 24512
rect 27556 24448 27564 24512
rect 27244 24447 27564 24448
rect 1744 23968 2064 23969
rect 1744 23904 1752 23968
rect 1816 23904 1832 23968
rect 1896 23904 1912 23968
rect 1976 23904 1992 23968
rect 2056 23904 2064 23968
rect 1744 23903 2064 23904
rect 4744 23968 5064 23969
rect 4744 23904 4752 23968
rect 4816 23904 4832 23968
rect 4896 23904 4912 23968
rect 4976 23904 4992 23968
rect 5056 23904 5064 23968
rect 4744 23903 5064 23904
rect 7744 23968 8064 23969
rect 7744 23904 7752 23968
rect 7816 23904 7832 23968
rect 7896 23904 7912 23968
rect 7976 23904 7992 23968
rect 8056 23904 8064 23968
rect 7744 23903 8064 23904
rect 10744 23968 11064 23969
rect 10744 23904 10752 23968
rect 10816 23904 10832 23968
rect 10896 23904 10912 23968
rect 10976 23904 10992 23968
rect 11056 23904 11064 23968
rect 10744 23903 11064 23904
rect 13744 23968 14064 23969
rect 13744 23904 13752 23968
rect 13816 23904 13832 23968
rect 13896 23904 13912 23968
rect 13976 23904 13992 23968
rect 14056 23904 14064 23968
rect 13744 23903 14064 23904
rect 16744 23968 17064 23969
rect 16744 23904 16752 23968
rect 16816 23904 16832 23968
rect 16896 23904 16912 23968
rect 16976 23904 16992 23968
rect 17056 23904 17064 23968
rect 16744 23903 17064 23904
rect 19744 23968 20064 23969
rect 19744 23904 19752 23968
rect 19816 23904 19832 23968
rect 19896 23904 19912 23968
rect 19976 23904 19992 23968
rect 20056 23904 20064 23968
rect 19744 23903 20064 23904
rect 22744 23968 23064 23969
rect 22744 23904 22752 23968
rect 22816 23904 22832 23968
rect 22896 23904 22912 23968
rect 22976 23904 22992 23968
rect 23056 23904 23064 23968
rect 22744 23903 23064 23904
rect 25744 23968 26064 23969
rect 25744 23904 25752 23968
rect 25816 23904 25832 23968
rect 25896 23904 25912 23968
rect 25976 23904 25992 23968
rect 26056 23904 26064 23968
rect 25744 23903 26064 23904
rect 3244 23424 3564 23425
rect 3244 23360 3252 23424
rect 3316 23360 3332 23424
rect 3396 23360 3412 23424
rect 3476 23360 3492 23424
rect 3556 23360 3564 23424
rect 3244 23359 3564 23360
rect 6244 23424 6564 23425
rect 6244 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6412 23424
rect 6476 23360 6492 23424
rect 6556 23360 6564 23424
rect 6244 23359 6564 23360
rect 9244 23424 9564 23425
rect 9244 23360 9252 23424
rect 9316 23360 9332 23424
rect 9396 23360 9412 23424
rect 9476 23360 9492 23424
rect 9556 23360 9564 23424
rect 9244 23359 9564 23360
rect 12244 23424 12564 23425
rect 12244 23360 12252 23424
rect 12316 23360 12332 23424
rect 12396 23360 12412 23424
rect 12476 23360 12492 23424
rect 12556 23360 12564 23424
rect 12244 23359 12564 23360
rect 15244 23424 15564 23425
rect 15244 23360 15252 23424
rect 15316 23360 15332 23424
rect 15396 23360 15412 23424
rect 15476 23360 15492 23424
rect 15556 23360 15564 23424
rect 15244 23359 15564 23360
rect 18244 23424 18564 23425
rect 18244 23360 18252 23424
rect 18316 23360 18332 23424
rect 18396 23360 18412 23424
rect 18476 23360 18492 23424
rect 18556 23360 18564 23424
rect 18244 23359 18564 23360
rect 21244 23424 21564 23425
rect 21244 23360 21252 23424
rect 21316 23360 21332 23424
rect 21396 23360 21412 23424
rect 21476 23360 21492 23424
rect 21556 23360 21564 23424
rect 21244 23359 21564 23360
rect 24244 23424 24564 23425
rect 24244 23360 24252 23424
rect 24316 23360 24332 23424
rect 24396 23360 24412 23424
rect 24476 23360 24492 23424
rect 24556 23360 24564 23424
rect 24244 23359 24564 23360
rect 27244 23424 27564 23425
rect 27244 23360 27252 23424
rect 27316 23360 27332 23424
rect 27396 23360 27412 23424
rect 27476 23360 27492 23424
rect 27556 23360 27564 23424
rect 27244 23359 27564 23360
rect 1744 22880 2064 22881
rect 1744 22816 1752 22880
rect 1816 22816 1832 22880
rect 1896 22816 1912 22880
rect 1976 22816 1992 22880
rect 2056 22816 2064 22880
rect 1744 22815 2064 22816
rect 4744 22880 5064 22881
rect 4744 22816 4752 22880
rect 4816 22816 4832 22880
rect 4896 22816 4912 22880
rect 4976 22816 4992 22880
rect 5056 22816 5064 22880
rect 4744 22815 5064 22816
rect 7744 22880 8064 22881
rect 7744 22816 7752 22880
rect 7816 22816 7832 22880
rect 7896 22816 7912 22880
rect 7976 22816 7992 22880
rect 8056 22816 8064 22880
rect 7744 22815 8064 22816
rect 10744 22880 11064 22881
rect 10744 22816 10752 22880
rect 10816 22816 10832 22880
rect 10896 22816 10912 22880
rect 10976 22816 10992 22880
rect 11056 22816 11064 22880
rect 10744 22815 11064 22816
rect 13744 22880 14064 22881
rect 13744 22816 13752 22880
rect 13816 22816 13832 22880
rect 13896 22816 13912 22880
rect 13976 22816 13992 22880
rect 14056 22816 14064 22880
rect 13744 22815 14064 22816
rect 16744 22880 17064 22881
rect 16744 22816 16752 22880
rect 16816 22816 16832 22880
rect 16896 22816 16912 22880
rect 16976 22816 16992 22880
rect 17056 22816 17064 22880
rect 16744 22815 17064 22816
rect 19744 22880 20064 22881
rect 19744 22816 19752 22880
rect 19816 22816 19832 22880
rect 19896 22816 19912 22880
rect 19976 22816 19992 22880
rect 20056 22816 20064 22880
rect 19744 22815 20064 22816
rect 22744 22880 23064 22881
rect 22744 22816 22752 22880
rect 22816 22816 22832 22880
rect 22896 22816 22912 22880
rect 22976 22816 22992 22880
rect 23056 22816 23064 22880
rect 22744 22815 23064 22816
rect 25744 22880 26064 22881
rect 25744 22816 25752 22880
rect 25816 22816 25832 22880
rect 25896 22816 25912 22880
rect 25976 22816 25992 22880
rect 26056 22816 26064 22880
rect 25744 22815 26064 22816
rect 3244 22336 3564 22337
rect 3244 22272 3252 22336
rect 3316 22272 3332 22336
rect 3396 22272 3412 22336
rect 3476 22272 3492 22336
rect 3556 22272 3564 22336
rect 3244 22271 3564 22272
rect 6244 22336 6564 22337
rect 6244 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6412 22336
rect 6476 22272 6492 22336
rect 6556 22272 6564 22336
rect 6244 22271 6564 22272
rect 9244 22336 9564 22337
rect 9244 22272 9252 22336
rect 9316 22272 9332 22336
rect 9396 22272 9412 22336
rect 9476 22272 9492 22336
rect 9556 22272 9564 22336
rect 9244 22271 9564 22272
rect 12244 22336 12564 22337
rect 12244 22272 12252 22336
rect 12316 22272 12332 22336
rect 12396 22272 12412 22336
rect 12476 22272 12492 22336
rect 12556 22272 12564 22336
rect 12244 22271 12564 22272
rect 15244 22336 15564 22337
rect 15244 22272 15252 22336
rect 15316 22272 15332 22336
rect 15396 22272 15412 22336
rect 15476 22272 15492 22336
rect 15556 22272 15564 22336
rect 15244 22271 15564 22272
rect 18244 22336 18564 22337
rect 18244 22272 18252 22336
rect 18316 22272 18332 22336
rect 18396 22272 18412 22336
rect 18476 22272 18492 22336
rect 18556 22272 18564 22336
rect 18244 22271 18564 22272
rect 21244 22336 21564 22337
rect 21244 22272 21252 22336
rect 21316 22272 21332 22336
rect 21396 22272 21412 22336
rect 21476 22272 21492 22336
rect 21556 22272 21564 22336
rect 21244 22271 21564 22272
rect 24244 22336 24564 22337
rect 24244 22272 24252 22336
rect 24316 22272 24332 22336
rect 24396 22272 24412 22336
rect 24476 22272 24492 22336
rect 24556 22272 24564 22336
rect 24244 22271 24564 22272
rect 27244 22336 27564 22337
rect 27244 22272 27252 22336
rect 27316 22272 27332 22336
rect 27396 22272 27412 22336
rect 27476 22272 27492 22336
rect 27556 22272 27564 22336
rect 27244 22271 27564 22272
rect 1744 21792 2064 21793
rect 1744 21728 1752 21792
rect 1816 21728 1832 21792
rect 1896 21728 1912 21792
rect 1976 21728 1992 21792
rect 2056 21728 2064 21792
rect 1744 21727 2064 21728
rect 4744 21792 5064 21793
rect 4744 21728 4752 21792
rect 4816 21728 4832 21792
rect 4896 21728 4912 21792
rect 4976 21728 4992 21792
rect 5056 21728 5064 21792
rect 4744 21727 5064 21728
rect 7744 21792 8064 21793
rect 7744 21728 7752 21792
rect 7816 21728 7832 21792
rect 7896 21728 7912 21792
rect 7976 21728 7992 21792
rect 8056 21728 8064 21792
rect 7744 21727 8064 21728
rect 10744 21792 11064 21793
rect 10744 21728 10752 21792
rect 10816 21728 10832 21792
rect 10896 21728 10912 21792
rect 10976 21728 10992 21792
rect 11056 21728 11064 21792
rect 10744 21727 11064 21728
rect 13744 21792 14064 21793
rect 13744 21728 13752 21792
rect 13816 21728 13832 21792
rect 13896 21728 13912 21792
rect 13976 21728 13992 21792
rect 14056 21728 14064 21792
rect 13744 21727 14064 21728
rect 16744 21792 17064 21793
rect 16744 21728 16752 21792
rect 16816 21728 16832 21792
rect 16896 21728 16912 21792
rect 16976 21728 16992 21792
rect 17056 21728 17064 21792
rect 16744 21727 17064 21728
rect 19744 21792 20064 21793
rect 19744 21728 19752 21792
rect 19816 21728 19832 21792
rect 19896 21728 19912 21792
rect 19976 21728 19992 21792
rect 20056 21728 20064 21792
rect 19744 21727 20064 21728
rect 22744 21792 23064 21793
rect 22744 21728 22752 21792
rect 22816 21728 22832 21792
rect 22896 21728 22912 21792
rect 22976 21728 22992 21792
rect 23056 21728 23064 21792
rect 22744 21727 23064 21728
rect 25744 21792 26064 21793
rect 25744 21728 25752 21792
rect 25816 21728 25832 21792
rect 25896 21728 25912 21792
rect 25976 21728 25992 21792
rect 26056 21728 26064 21792
rect 25744 21727 26064 21728
rect 3244 21248 3564 21249
rect 3244 21184 3252 21248
rect 3316 21184 3332 21248
rect 3396 21184 3412 21248
rect 3476 21184 3492 21248
rect 3556 21184 3564 21248
rect 3244 21183 3564 21184
rect 6244 21248 6564 21249
rect 6244 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6412 21248
rect 6476 21184 6492 21248
rect 6556 21184 6564 21248
rect 6244 21183 6564 21184
rect 9244 21248 9564 21249
rect 9244 21184 9252 21248
rect 9316 21184 9332 21248
rect 9396 21184 9412 21248
rect 9476 21184 9492 21248
rect 9556 21184 9564 21248
rect 9244 21183 9564 21184
rect 12244 21248 12564 21249
rect 12244 21184 12252 21248
rect 12316 21184 12332 21248
rect 12396 21184 12412 21248
rect 12476 21184 12492 21248
rect 12556 21184 12564 21248
rect 12244 21183 12564 21184
rect 15244 21248 15564 21249
rect 15244 21184 15252 21248
rect 15316 21184 15332 21248
rect 15396 21184 15412 21248
rect 15476 21184 15492 21248
rect 15556 21184 15564 21248
rect 15244 21183 15564 21184
rect 18244 21248 18564 21249
rect 18244 21184 18252 21248
rect 18316 21184 18332 21248
rect 18396 21184 18412 21248
rect 18476 21184 18492 21248
rect 18556 21184 18564 21248
rect 18244 21183 18564 21184
rect 21244 21248 21564 21249
rect 21244 21184 21252 21248
rect 21316 21184 21332 21248
rect 21396 21184 21412 21248
rect 21476 21184 21492 21248
rect 21556 21184 21564 21248
rect 21244 21183 21564 21184
rect 24244 21248 24564 21249
rect 24244 21184 24252 21248
rect 24316 21184 24332 21248
rect 24396 21184 24412 21248
rect 24476 21184 24492 21248
rect 24556 21184 24564 21248
rect 24244 21183 24564 21184
rect 27244 21248 27564 21249
rect 27244 21184 27252 21248
rect 27316 21184 27332 21248
rect 27396 21184 27412 21248
rect 27476 21184 27492 21248
rect 27556 21184 27564 21248
rect 27244 21183 27564 21184
rect 1744 20704 2064 20705
rect 1744 20640 1752 20704
rect 1816 20640 1832 20704
rect 1896 20640 1912 20704
rect 1976 20640 1992 20704
rect 2056 20640 2064 20704
rect 1744 20639 2064 20640
rect 4744 20704 5064 20705
rect 4744 20640 4752 20704
rect 4816 20640 4832 20704
rect 4896 20640 4912 20704
rect 4976 20640 4992 20704
rect 5056 20640 5064 20704
rect 4744 20639 5064 20640
rect 7744 20704 8064 20705
rect 7744 20640 7752 20704
rect 7816 20640 7832 20704
rect 7896 20640 7912 20704
rect 7976 20640 7992 20704
rect 8056 20640 8064 20704
rect 7744 20639 8064 20640
rect 10744 20704 11064 20705
rect 10744 20640 10752 20704
rect 10816 20640 10832 20704
rect 10896 20640 10912 20704
rect 10976 20640 10992 20704
rect 11056 20640 11064 20704
rect 10744 20639 11064 20640
rect 13744 20704 14064 20705
rect 13744 20640 13752 20704
rect 13816 20640 13832 20704
rect 13896 20640 13912 20704
rect 13976 20640 13992 20704
rect 14056 20640 14064 20704
rect 13744 20639 14064 20640
rect 16744 20704 17064 20705
rect 16744 20640 16752 20704
rect 16816 20640 16832 20704
rect 16896 20640 16912 20704
rect 16976 20640 16992 20704
rect 17056 20640 17064 20704
rect 16744 20639 17064 20640
rect 19744 20704 20064 20705
rect 19744 20640 19752 20704
rect 19816 20640 19832 20704
rect 19896 20640 19912 20704
rect 19976 20640 19992 20704
rect 20056 20640 20064 20704
rect 19744 20639 20064 20640
rect 22744 20704 23064 20705
rect 22744 20640 22752 20704
rect 22816 20640 22832 20704
rect 22896 20640 22912 20704
rect 22976 20640 22992 20704
rect 23056 20640 23064 20704
rect 22744 20639 23064 20640
rect 25744 20704 26064 20705
rect 25744 20640 25752 20704
rect 25816 20640 25832 20704
rect 25896 20640 25912 20704
rect 25976 20640 25992 20704
rect 26056 20640 26064 20704
rect 25744 20639 26064 20640
rect 3244 20160 3564 20161
rect 3244 20096 3252 20160
rect 3316 20096 3332 20160
rect 3396 20096 3412 20160
rect 3476 20096 3492 20160
rect 3556 20096 3564 20160
rect 3244 20095 3564 20096
rect 6244 20160 6564 20161
rect 6244 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6412 20160
rect 6476 20096 6492 20160
rect 6556 20096 6564 20160
rect 6244 20095 6564 20096
rect 9244 20160 9564 20161
rect 9244 20096 9252 20160
rect 9316 20096 9332 20160
rect 9396 20096 9412 20160
rect 9476 20096 9492 20160
rect 9556 20096 9564 20160
rect 9244 20095 9564 20096
rect 12244 20160 12564 20161
rect 12244 20096 12252 20160
rect 12316 20096 12332 20160
rect 12396 20096 12412 20160
rect 12476 20096 12492 20160
rect 12556 20096 12564 20160
rect 12244 20095 12564 20096
rect 15244 20160 15564 20161
rect 15244 20096 15252 20160
rect 15316 20096 15332 20160
rect 15396 20096 15412 20160
rect 15476 20096 15492 20160
rect 15556 20096 15564 20160
rect 15244 20095 15564 20096
rect 18244 20160 18564 20161
rect 18244 20096 18252 20160
rect 18316 20096 18332 20160
rect 18396 20096 18412 20160
rect 18476 20096 18492 20160
rect 18556 20096 18564 20160
rect 18244 20095 18564 20096
rect 21244 20160 21564 20161
rect 21244 20096 21252 20160
rect 21316 20096 21332 20160
rect 21396 20096 21412 20160
rect 21476 20096 21492 20160
rect 21556 20096 21564 20160
rect 21244 20095 21564 20096
rect 24244 20160 24564 20161
rect 24244 20096 24252 20160
rect 24316 20096 24332 20160
rect 24396 20096 24412 20160
rect 24476 20096 24492 20160
rect 24556 20096 24564 20160
rect 24244 20095 24564 20096
rect 27244 20160 27564 20161
rect 27244 20096 27252 20160
rect 27316 20096 27332 20160
rect 27396 20096 27412 20160
rect 27476 20096 27492 20160
rect 27556 20096 27564 20160
rect 27244 20095 27564 20096
rect 1744 19616 2064 19617
rect 1744 19552 1752 19616
rect 1816 19552 1832 19616
rect 1896 19552 1912 19616
rect 1976 19552 1992 19616
rect 2056 19552 2064 19616
rect 1744 19551 2064 19552
rect 4744 19616 5064 19617
rect 4744 19552 4752 19616
rect 4816 19552 4832 19616
rect 4896 19552 4912 19616
rect 4976 19552 4992 19616
rect 5056 19552 5064 19616
rect 4744 19551 5064 19552
rect 7744 19616 8064 19617
rect 7744 19552 7752 19616
rect 7816 19552 7832 19616
rect 7896 19552 7912 19616
rect 7976 19552 7992 19616
rect 8056 19552 8064 19616
rect 7744 19551 8064 19552
rect 10744 19616 11064 19617
rect 10744 19552 10752 19616
rect 10816 19552 10832 19616
rect 10896 19552 10912 19616
rect 10976 19552 10992 19616
rect 11056 19552 11064 19616
rect 10744 19551 11064 19552
rect 13744 19616 14064 19617
rect 13744 19552 13752 19616
rect 13816 19552 13832 19616
rect 13896 19552 13912 19616
rect 13976 19552 13992 19616
rect 14056 19552 14064 19616
rect 13744 19551 14064 19552
rect 16744 19616 17064 19617
rect 16744 19552 16752 19616
rect 16816 19552 16832 19616
rect 16896 19552 16912 19616
rect 16976 19552 16992 19616
rect 17056 19552 17064 19616
rect 16744 19551 17064 19552
rect 19744 19616 20064 19617
rect 19744 19552 19752 19616
rect 19816 19552 19832 19616
rect 19896 19552 19912 19616
rect 19976 19552 19992 19616
rect 20056 19552 20064 19616
rect 19744 19551 20064 19552
rect 22744 19616 23064 19617
rect 22744 19552 22752 19616
rect 22816 19552 22832 19616
rect 22896 19552 22912 19616
rect 22976 19552 22992 19616
rect 23056 19552 23064 19616
rect 22744 19551 23064 19552
rect 25744 19616 26064 19617
rect 25744 19552 25752 19616
rect 25816 19552 25832 19616
rect 25896 19552 25912 19616
rect 25976 19552 25992 19616
rect 26056 19552 26064 19616
rect 25744 19551 26064 19552
rect 3244 19072 3564 19073
rect 3244 19008 3252 19072
rect 3316 19008 3332 19072
rect 3396 19008 3412 19072
rect 3476 19008 3492 19072
rect 3556 19008 3564 19072
rect 3244 19007 3564 19008
rect 6244 19072 6564 19073
rect 6244 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6412 19072
rect 6476 19008 6492 19072
rect 6556 19008 6564 19072
rect 6244 19007 6564 19008
rect 9244 19072 9564 19073
rect 9244 19008 9252 19072
rect 9316 19008 9332 19072
rect 9396 19008 9412 19072
rect 9476 19008 9492 19072
rect 9556 19008 9564 19072
rect 9244 19007 9564 19008
rect 12244 19072 12564 19073
rect 12244 19008 12252 19072
rect 12316 19008 12332 19072
rect 12396 19008 12412 19072
rect 12476 19008 12492 19072
rect 12556 19008 12564 19072
rect 12244 19007 12564 19008
rect 15244 19072 15564 19073
rect 15244 19008 15252 19072
rect 15316 19008 15332 19072
rect 15396 19008 15412 19072
rect 15476 19008 15492 19072
rect 15556 19008 15564 19072
rect 15244 19007 15564 19008
rect 18244 19072 18564 19073
rect 18244 19008 18252 19072
rect 18316 19008 18332 19072
rect 18396 19008 18412 19072
rect 18476 19008 18492 19072
rect 18556 19008 18564 19072
rect 18244 19007 18564 19008
rect 21244 19072 21564 19073
rect 21244 19008 21252 19072
rect 21316 19008 21332 19072
rect 21396 19008 21412 19072
rect 21476 19008 21492 19072
rect 21556 19008 21564 19072
rect 21244 19007 21564 19008
rect 24244 19072 24564 19073
rect 24244 19008 24252 19072
rect 24316 19008 24332 19072
rect 24396 19008 24412 19072
rect 24476 19008 24492 19072
rect 24556 19008 24564 19072
rect 24244 19007 24564 19008
rect 27244 19072 27564 19073
rect 27244 19008 27252 19072
rect 27316 19008 27332 19072
rect 27396 19008 27412 19072
rect 27476 19008 27492 19072
rect 27556 19008 27564 19072
rect 27244 19007 27564 19008
rect 1744 18528 2064 18529
rect 1744 18464 1752 18528
rect 1816 18464 1832 18528
rect 1896 18464 1912 18528
rect 1976 18464 1992 18528
rect 2056 18464 2064 18528
rect 1744 18463 2064 18464
rect 4744 18528 5064 18529
rect 4744 18464 4752 18528
rect 4816 18464 4832 18528
rect 4896 18464 4912 18528
rect 4976 18464 4992 18528
rect 5056 18464 5064 18528
rect 4744 18463 5064 18464
rect 7744 18528 8064 18529
rect 7744 18464 7752 18528
rect 7816 18464 7832 18528
rect 7896 18464 7912 18528
rect 7976 18464 7992 18528
rect 8056 18464 8064 18528
rect 7744 18463 8064 18464
rect 10744 18528 11064 18529
rect 10744 18464 10752 18528
rect 10816 18464 10832 18528
rect 10896 18464 10912 18528
rect 10976 18464 10992 18528
rect 11056 18464 11064 18528
rect 10744 18463 11064 18464
rect 13744 18528 14064 18529
rect 13744 18464 13752 18528
rect 13816 18464 13832 18528
rect 13896 18464 13912 18528
rect 13976 18464 13992 18528
rect 14056 18464 14064 18528
rect 13744 18463 14064 18464
rect 16744 18528 17064 18529
rect 16744 18464 16752 18528
rect 16816 18464 16832 18528
rect 16896 18464 16912 18528
rect 16976 18464 16992 18528
rect 17056 18464 17064 18528
rect 16744 18463 17064 18464
rect 19744 18528 20064 18529
rect 19744 18464 19752 18528
rect 19816 18464 19832 18528
rect 19896 18464 19912 18528
rect 19976 18464 19992 18528
rect 20056 18464 20064 18528
rect 19744 18463 20064 18464
rect 22744 18528 23064 18529
rect 22744 18464 22752 18528
rect 22816 18464 22832 18528
rect 22896 18464 22912 18528
rect 22976 18464 22992 18528
rect 23056 18464 23064 18528
rect 22744 18463 23064 18464
rect 25744 18528 26064 18529
rect 25744 18464 25752 18528
rect 25816 18464 25832 18528
rect 25896 18464 25912 18528
rect 25976 18464 25992 18528
rect 26056 18464 26064 18528
rect 25744 18463 26064 18464
rect 3244 17984 3564 17985
rect 3244 17920 3252 17984
rect 3316 17920 3332 17984
rect 3396 17920 3412 17984
rect 3476 17920 3492 17984
rect 3556 17920 3564 17984
rect 3244 17919 3564 17920
rect 6244 17984 6564 17985
rect 6244 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6412 17984
rect 6476 17920 6492 17984
rect 6556 17920 6564 17984
rect 6244 17919 6564 17920
rect 9244 17984 9564 17985
rect 9244 17920 9252 17984
rect 9316 17920 9332 17984
rect 9396 17920 9412 17984
rect 9476 17920 9492 17984
rect 9556 17920 9564 17984
rect 9244 17919 9564 17920
rect 12244 17984 12564 17985
rect 12244 17920 12252 17984
rect 12316 17920 12332 17984
rect 12396 17920 12412 17984
rect 12476 17920 12492 17984
rect 12556 17920 12564 17984
rect 12244 17919 12564 17920
rect 15244 17984 15564 17985
rect 15244 17920 15252 17984
rect 15316 17920 15332 17984
rect 15396 17920 15412 17984
rect 15476 17920 15492 17984
rect 15556 17920 15564 17984
rect 15244 17919 15564 17920
rect 18244 17984 18564 17985
rect 18244 17920 18252 17984
rect 18316 17920 18332 17984
rect 18396 17920 18412 17984
rect 18476 17920 18492 17984
rect 18556 17920 18564 17984
rect 18244 17919 18564 17920
rect 21244 17984 21564 17985
rect 21244 17920 21252 17984
rect 21316 17920 21332 17984
rect 21396 17920 21412 17984
rect 21476 17920 21492 17984
rect 21556 17920 21564 17984
rect 21244 17919 21564 17920
rect 24244 17984 24564 17985
rect 24244 17920 24252 17984
rect 24316 17920 24332 17984
rect 24396 17920 24412 17984
rect 24476 17920 24492 17984
rect 24556 17920 24564 17984
rect 24244 17919 24564 17920
rect 27244 17984 27564 17985
rect 27244 17920 27252 17984
rect 27316 17920 27332 17984
rect 27396 17920 27412 17984
rect 27476 17920 27492 17984
rect 27556 17920 27564 17984
rect 27244 17919 27564 17920
rect 1744 17440 2064 17441
rect 1744 17376 1752 17440
rect 1816 17376 1832 17440
rect 1896 17376 1912 17440
rect 1976 17376 1992 17440
rect 2056 17376 2064 17440
rect 1744 17375 2064 17376
rect 4744 17440 5064 17441
rect 4744 17376 4752 17440
rect 4816 17376 4832 17440
rect 4896 17376 4912 17440
rect 4976 17376 4992 17440
rect 5056 17376 5064 17440
rect 4744 17375 5064 17376
rect 7744 17440 8064 17441
rect 7744 17376 7752 17440
rect 7816 17376 7832 17440
rect 7896 17376 7912 17440
rect 7976 17376 7992 17440
rect 8056 17376 8064 17440
rect 7744 17375 8064 17376
rect 10744 17440 11064 17441
rect 10744 17376 10752 17440
rect 10816 17376 10832 17440
rect 10896 17376 10912 17440
rect 10976 17376 10992 17440
rect 11056 17376 11064 17440
rect 10744 17375 11064 17376
rect 13744 17440 14064 17441
rect 13744 17376 13752 17440
rect 13816 17376 13832 17440
rect 13896 17376 13912 17440
rect 13976 17376 13992 17440
rect 14056 17376 14064 17440
rect 13744 17375 14064 17376
rect 16744 17440 17064 17441
rect 16744 17376 16752 17440
rect 16816 17376 16832 17440
rect 16896 17376 16912 17440
rect 16976 17376 16992 17440
rect 17056 17376 17064 17440
rect 16744 17375 17064 17376
rect 19744 17440 20064 17441
rect 19744 17376 19752 17440
rect 19816 17376 19832 17440
rect 19896 17376 19912 17440
rect 19976 17376 19992 17440
rect 20056 17376 20064 17440
rect 19744 17375 20064 17376
rect 22744 17440 23064 17441
rect 22744 17376 22752 17440
rect 22816 17376 22832 17440
rect 22896 17376 22912 17440
rect 22976 17376 22992 17440
rect 23056 17376 23064 17440
rect 22744 17375 23064 17376
rect 25744 17440 26064 17441
rect 25744 17376 25752 17440
rect 25816 17376 25832 17440
rect 25896 17376 25912 17440
rect 25976 17376 25992 17440
rect 26056 17376 26064 17440
rect 25744 17375 26064 17376
rect 3244 16896 3564 16897
rect 3244 16832 3252 16896
rect 3316 16832 3332 16896
rect 3396 16832 3412 16896
rect 3476 16832 3492 16896
rect 3556 16832 3564 16896
rect 3244 16831 3564 16832
rect 6244 16896 6564 16897
rect 6244 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6412 16896
rect 6476 16832 6492 16896
rect 6556 16832 6564 16896
rect 6244 16831 6564 16832
rect 9244 16896 9564 16897
rect 9244 16832 9252 16896
rect 9316 16832 9332 16896
rect 9396 16832 9412 16896
rect 9476 16832 9492 16896
rect 9556 16832 9564 16896
rect 9244 16831 9564 16832
rect 12244 16896 12564 16897
rect 12244 16832 12252 16896
rect 12316 16832 12332 16896
rect 12396 16832 12412 16896
rect 12476 16832 12492 16896
rect 12556 16832 12564 16896
rect 12244 16831 12564 16832
rect 15244 16896 15564 16897
rect 15244 16832 15252 16896
rect 15316 16832 15332 16896
rect 15396 16832 15412 16896
rect 15476 16832 15492 16896
rect 15556 16832 15564 16896
rect 15244 16831 15564 16832
rect 18244 16896 18564 16897
rect 18244 16832 18252 16896
rect 18316 16832 18332 16896
rect 18396 16832 18412 16896
rect 18476 16832 18492 16896
rect 18556 16832 18564 16896
rect 18244 16831 18564 16832
rect 21244 16896 21564 16897
rect 21244 16832 21252 16896
rect 21316 16832 21332 16896
rect 21396 16832 21412 16896
rect 21476 16832 21492 16896
rect 21556 16832 21564 16896
rect 21244 16831 21564 16832
rect 24244 16896 24564 16897
rect 24244 16832 24252 16896
rect 24316 16832 24332 16896
rect 24396 16832 24412 16896
rect 24476 16832 24492 16896
rect 24556 16832 24564 16896
rect 24244 16831 24564 16832
rect 27244 16896 27564 16897
rect 27244 16832 27252 16896
rect 27316 16832 27332 16896
rect 27396 16832 27412 16896
rect 27476 16832 27492 16896
rect 27556 16832 27564 16896
rect 27244 16831 27564 16832
rect 1744 16352 2064 16353
rect 1744 16288 1752 16352
rect 1816 16288 1832 16352
rect 1896 16288 1912 16352
rect 1976 16288 1992 16352
rect 2056 16288 2064 16352
rect 1744 16287 2064 16288
rect 4744 16352 5064 16353
rect 4744 16288 4752 16352
rect 4816 16288 4832 16352
rect 4896 16288 4912 16352
rect 4976 16288 4992 16352
rect 5056 16288 5064 16352
rect 4744 16287 5064 16288
rect 7744 16352 8064 16353
rect 7744 16288 7752 16352
rect 7816 16288 7832 16352
rect 7896 16288 7912 16352
rect 7976 16288 7992 16352
rect 8056 16288 8064 16352
rect 7744 16287 8064 16288
rect 10744 16352 11064 16353
rect 10744 16288 10752 16352
rect 10816 16288 10832 16352
rect 10896 16288 10912 16352
rect 10976 16288 10992 16352
rect 11056 16288 11064 16352
rect 10744 16287 11064 16288
rect 13744 16352 14064 16353
rect 13744 16288 13752 16352
rect 13816 16288 13832 16352
rect 13896 16288 13912 16352
rect 13976 16288 13992 16352
rect 14056 16288 14064 16352
rect 13744 16287 14064 16288
rect 16744 16352 17064 16353
rect 16744 16288 16752 16352
rect 16816 16288 16832 16352
rect 16896 16288 16912 16352
rect 16976 16288 16992 16352
rect 17056 16288 17064 16352
rect 16744 16287 17064 16288
rect 19744 16352 20064 16353
rect 19744 16288 19752 16352
rect 19816 16288 19832 16352
rect 19896 16288 19912 16352
rect 19976 16288 19992 16352
rect 20056 16288 20064 16352
rect 19744 16287 20064 16288
rect 22744 16352 23064 16353
rect 22744 16288 22752 16352
rect 22816 16288 22832 16352
rect 22896 16288 22912 16352
rect 22976 16288 22992 16352
rect 23056 16288 23064 16352
rect 22744 16287 23064 16288
rect 25744 16352 26064 16353
rect 25744 16288 25752 16352
rect 25816 16288 25832 16352
rect 25896 16288 25912 16352
rect 25976 16288 25992 16352
rect 26056 16288 26064 16352
rect 25744 16287 26064 16288
rect 3244 15808 3564 15809
rect 3244 15744 3252 15808
rect 3316 15744 3332 15808
rect 3396 15744 3412 15808
rect 3476 15744 3492 15808
rect 3556 15744 3564 15808
rect 3244 15743 3564 15744
rect 6244 15808 6564 15809
rect 6244 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6412 15808
rect 6476 15744 6492 15808
rect 6556 15744 6564 15808
rect 6244 15743 6564 15744
rect 9244 15808 9564 15809
rect 9244 15744 9252 15808
rect 9316 15744 9332 15808
rect 9396 15744 9412 15808
rect 9476 15744 9492 15808
rect 9556 15744 9564 15808
rect 9244 15743 9564 15744
rect 12244 15808 12564 15809
rect 12244 15744 12252 15808
rect 12316 15744 12332 15808
rect 12396 15744 12412 15808
rect 12476 15744 12492 15808
rect 12556 15744 12564 15808
rect 12244 15743 12564 15744
rect 15244 15808 15564 15809
rect 15244 15744 15252 15808
rect 15316 15744 15332 15808
rect 15396 15744 15412 15808
rect 15476 15744 15492 15808
rect 15556 15744 15564 15808
rect 15244 15743 15564 15744
rect 18244 15808 18564 15809
rect 18244 15744 18252 15808
rect 18316 15744 18332 15808
rect 18396 15744 18412 15808
rect 18476 15744 18492 15808
rect 18556 15744 18564 15808
rect 18244 15743 18564 15744
rect 21244 15808 21564 15809
rect 21244 15744 21252 15808
rect 21316 15744 21332 15808
rect 21396 15744 21412 15808
rect 21476 15744 21492 15808
rect 21556 15744 21564 15808
rect 21244 15743 21564 15744
rect 24244 15808 24564 15809
rect 24244 15744 24252 15808
rect 24316 15744 24332 15808
rect 24396 15744 24412 15808
rect 24476 15744 24492 15808
rect 24556 15744 24564 15808
rect 24244 15743 24564 15744
rect 27244 15808 27564 15809
rect 27244 15744 27252 15808
rect 27316 15744 27332 15808
rect 27396 15744 27412 15808
rect 27476 15744 27492 15808
rect 27556 15744 27564 15808
rect 27244 15743 27564 15744
rect 1744 15264 2064 15265
rect 1744 15200 1752 15264
rect 1816 15200 1832 15264
rect 1896 15200 1912 15264
rect 1976 15200 1992 15264
rect 2056 15200 2064 15264
rect 1744 15199 2064 15200
rect 4744 15264 5064 15265
rect 4744 15200 4752 15264
rect 4816 15200 4832 15264
rect 4896 15200 4912 15264
rect 4976 15200 4992 15264
rect 5056 15200 5064 15264
rect 4744 15199 5064 15200
rect 7744 15264 8064 15265
rect 7744 15200 7752 15264
rect 7816 15200 7832 15264
rect 7896 15200 7912 15264
rect 7976 15200 7992 15264
rect 8056 15200 8064 15264
rect 7744 15199 8064 15200
rect 10744 15264 11064 15265
rect 10744 15200 10752 15264
rect 10816 15200 10832 15264
rect 10896 15200 10912 15264
rect 10976 15200 10992 15264
rect 11056 15200 11064 15264
rect 10744 15199 11064 15200
rect 13744 15264 14064 15265
rect 13744 15200 13752 15264
rect 13816 15200 13832 15264
rect 13896 15200 13912 15264
rect 13976 15200 13992 15264
rect 14056 15200 14064 15264
rect 13744 15199 14064 15200
rect 16744 15264 17064 15265
rect 16744 15200 16752 15264
rect 16816 15200 16832 15264
rect 16896 15200 16912 15264
rect 16976 15200 16992 15264
rect 17056 15200 17064 15264
rect 16744 15199 17064 15200
rect 19744 15264 20064 15265
rect 19744 15200 19752 15264
rect 19816 15200 19832 15264
rect 19896 15200 19912 15264
rect 19976 15200 19992 15264
rect 20056 15200 20064 15264
rect 19744 15199 20064 15200
rect 22744 15264 23064 15265
rect 22744 15200 22752 15264
rect 22816 15200 22832 15264
rect 22896 15200 22912 15264
rect 22976 15200 22992 15264
rect 23056 15200 23064 15264
rect 22744 15199 23064 15200
rect 25744 15264 26064 15265
rect 25744 15200 25752 15264
rect 25816 15200 25832 15264
rect 25896 15200 25912 15264
rect 25976 15200 25992 15264
rect 26056 15200 26064 15264
rect 25744 15199 26064 15200
rect 3244 14720 3564 14721
rect 3244 14656 3252 14720
rect 3316 14656 3332 14720
rect 3396 14656 3412 14720
rect 3476 14656 3492 14720
rect 3556 14656 3564 14720
rect 3244 14655 3564 14656
rect 6244 14720 6564 14721
rect 6244 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6412 14720
rect 6476 14656 6492 14720
rect 6556 14656 6564 14720
rect 6244 14655 6564 14656
rect 9244 14720 9564 14721
rect 9244 14656 9252 14720
rect 9316 14656 9332 14720
rect 9396 14656 9412 14720
rect 9476 14656 9492 14720
rect 9556 14656 9564 14720
rect 9244 14655 9564 14656
rect 12244 14720 12564 14721
rect 12244 14656 12252 14720
rect 12316 14656 12332 14720
rect 12396 14656 12412 14720
rect 12476 14656 12492 14720
rect 12556 14656 12564 14720
rect 12244 14655 12564 14656
rect 15244 14720 15564 14721
rect 15244 14656 15252 14720
rect 15316 14656 15332 14720
rect 15396 14656 15412 14720
rect 15476 14656 15492 14720
rect 15556 14656 15564 14720
rect 15244 14655 15564 14656
rect 18244 14720 18564 14721
rect 18244 14656 18252 14720
rect 18316 14656 18332 14720
rect 18396 14656 18412 14720
rect 18476 14656 18492 14720
rect 18556 14656 18564 14720
rect 18244 14655 18564 14656
rect 21244 14720 21564 14721
rect 21244 14656 21252 14720
rect 21316 14656 21332 14720
rect 21396 14656 21412 14720
rect 21476 14656 21492 14720
rect 21556 14656 21564 14720
rect 21244 14655 21564 14656
rect 24244 14720 24564 14721
rect 24244 14656 24252 14720
rect 24316 14656 24332 14720
rect 24396 14656 24412 14720
rect 24476 14656 24492 14720
rect 24556 14656 24564 14720
rect 24244 14655 24564 14656
rect 27244 14720 27564 14721
rect 27244 14656 27252 14720
rect 27316 14656 27332 14720
rect 27396 14656 27412 14720
rect 27476 14656 27492 14720
rect 27556 14656 27564 14720
rect 27244 14655 27564 14656
rect 14273 14514 14339 14517
rect 19374 14514 19380 14516
rect 14273 14512 19380 14514
rect 14273 14456 14278 14512
rect 14334 14456 19380 14512
rect 14273 14454 19380 14456
rect 14273 14451 14339 14454
rect 19374 14452 19380 14454
rect 19444 14514 19450 14516
rect 21633 14514 21699 14517
rect 19444 14512 21699 14514
rect 19444 14456 21638 14512
rect 21694 14456 21699 14512
rect 19444 14454 21699 14456
rect 19444 14452 19450 14454
rect 21633 14451 21699 14454
rect 1744 14176 2064 14177
rect 1744 14112 1752 14176
rect 1816 14112 1832 14176
rect 1896 14112 1912 14176
rect 1976 14112 1992 14176
rect 2056 14112 2064 14176
rect 1744 14111 2064 14112
rect 4744 14176 5064 14177
rect 4744 14112 4752 14176
rect 4816 14112 4832 14176
rect 4896 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5064 14176
rect 4744 14111 5064 14112
rect 7744 14176 8064 14177
rect 7744 14112 7752 14176
rect 7816 14112 7832 14176
rect 7896 14112 7912 14176
rect 7976 14112 7992 14176
rect 8056 14112 8064 14176
rect 7744 14111 8064 14112
rect 10744 14176 11064 14177
rect 10744 14112 10752 14176
rect 10816 14112 10832 14176
rect 10896 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11064 14176
rect 10744 14111 11064 14112
rect 13744 14176 14064 14177
rect 13744 14112 13752 14176
rect 13816 14112 13832 14176
rect 13896 14112 13912 14176
rect 13976 14112 13992 14176
rect 14056 14112 14064 14176
rect 13744 14111 14064 14112
rect 16744 14176 17064 14177
rect 16744 14112 16752 14176
rect 16816 14112 16832 14176
rect 16896 14112 16912 14176
rect 16976 14112 16992 14176
rect 17056 14112 17064 14176
rect 16744 14111 17064 14112
rect 19744 14176 20064 14177
rect 19744 14112 19752 14176
rect 19816 14112 19832 14176
rect 19896 14112 19912 14176
rect 19976 14112 19992 14176
rect 20056 14112 20064 14176
rect 19744 14111 20064 14112
rect 22744 14176 23064 14177
rect 22744 14112 22752 14176
rect 22816 14112 22832 14176
rect 22896 14112 22912 14176
rect 22976 14112 22992 14176
rect 23056 14112 23064 14176
rect 22744 14111 23064 14112
rect 25744 14176 26064 14177
rect 25744 14112 25752 14176
rect 25816 14112 25832 14176
rect 25896 14112 25912 14176
rect 25976 14112 25992 14176
rect 26056 14112 26064 14176
rect 25744 14111 26064 14112
rect 8477 13970 8543 13973
rect 14089 13970 14155 13973
rect 8477 13968 14155 13970
rect 8477 13912 8482 13968
rect 8538 13912 14094 13968
rect 14150 13912 14155 13968
rect 8477 13910 14155 13912
rect 8477 13907 8543 13910
rect 14089 13907 14155 13910
rect 0 13696 800 13728
rect 0 13640 110 13696
rect 166 13640 800 13696
rect 0 13608 800 13640
rect 3244 13632 3564 13633
rect 3244 13568 3252 13632
rect 3316 13568 3332 13632
rect 3396 13568 3412 13632
rect 3476 13568 3492 13632
rect 3556 13568 3564 13632
rect 3244 13567 3564 13568
rect 6244 13632 6564 13633
rect 6244 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6412 13632
rect 6476 13568 6492 13632
rect 6556 13568 6564 13632
rect 6244 13567 6564 13568
rect 9244 13632 9564 13633
rect 9244 13568 9252 13632
rect 9316 13568 9332 13632
rect 9396 13568 9412 13632
rect 9476 13568 9492 13632
rect 9556 13568 9564 13632
rect 9244 13567 9564 13568
rect 12244 13632 12564 13633
rect 12244 13568 12252 13632
rect 12316 13568 12332 13632
rect 12396 13568 12412 13632
rect 12476 13568 12492 13632
rect 12556 13568 12564 13632
rect 12244 13567 12564 13568
rect 15244 13632 15564 13633
rect 15244 13568 15252 13632
rect 15316 13568 15332 13632
rect 15396 13568 15412 13632
rect 15476 13568 15492 13632
rect 15556 13568 15564 13632
rect 15244 13567 15564 13568
rect 18244 13632 18564 13633
rect 18244 13568 18252 13632
rect 18316 13568 18332 13632
rect 18396 13568 18412 13632
rect 18476 13568 18492 13632
rect 18556 13568 18564 13632
rect 18244 13567 18564 13568
rect 21244 13632 21564 13633
rect 21244 13568 21252 13632
rect 21316 13568 21332 13632
rect 21396 13568 21412 13632
rect 21476 13568 21492 13632
rect 21556 13568 21564 13632
rect 21244 13567 21564 13568
rect 24244 13632 24564 13633
rect 24244 13568 24252 13632
rect 24316 13568 24332 13632
rect 24396 13568 24412 13632
rect 24476 13568 24492 13632
rect 24556 13568 24564 13632
rect 24244 13567 24564 13568
rect 27244 13632 27564 13633
rect 27244 13568 27252 13632
rect 27316 13568 27332 13632
rect 27396 13568 27412 13632
rect 27476 13568 27492 13632
rect 27556 13568 27564 13632
rect 27244 13567 27564 13568
rect 1744 13088 2064 13089
rect 1744 13024 1752 13088
rect 1816 13024 1832 13088
rect 1896 13024 1912 13088
rect 1976 13024 1992 13088
rect 2056 13024 2064 13088
rect 1744 13023 2064 13024
rect 4744 13088 5064 13089
rect 4744 13024 4752 13088
rect 4816 13024 4832 13088
rect 4896 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5064 13088
rect 4744 13023 5064 13024
rect 7744 13088 8064 13089
rect 7744 13024 7752 13088
rect 7816 13024 7832 13088
rect 7896 13024 7912 13088
rect 7976 13024 7992 13088
rect 8056 13024 8064 13088
rect 7744 13023 8064 13024
rect 10744 13088 11064 13089
rect 10744 13024 10752 13088
rect 10816 13024 10832 13088
rect 10896 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11064 13088
rect 10744 13023 11064 13024
rect 13744 13088 14064 13089
rect 13744 13024 13752 13088
rect 13816 13024 13832 13088
rect 13896 13024 13912 13088
rect 13976 13024 13992 13088
rect 14056 13024 14064 13088
rect 13744 13023 14064 13024
rect 16744 13088 17064 13089
rect 16744 13024 16752 13088
rect 16816 13024 16832 13088
rect 16896 13024 16912 13088
rect 16976 13024 16992 13088
rect 17056 13024 17064 13088
rect 16744 13023 17064 13024
rect 19744 13088 20064 13089
rect 19744 13024 19752 13088
rect 19816 13024 19832 13088
rect 19896 13024 19912 13088
rect 19976 13024 19992 13088
rect 20056 13024 20064 13088
rect 19744 13023 20064 13024
rect 22744 13088 23064 13089
rect 22744 13024 22752 13088
rect 22816 13024 22832 13088
rect 22896 13024 22912 13088
rect 22976 13024 22992 13088
rect 23056 13024 23064 13088
rect 22744 13023 23064 13024
rect 25744 13088 26064 13089
rect 25744 13024 25752 13088
rect 25816 13024 25832 13088
rect 25896 13024 25912 13088
rect 25976 13024 25992 13088
rect 26056 13024 26064 13088
rect 25744 13023 26064 13024
rect 105 12746 171 12749
rect 23197 12746 23263 12749
rect 105 12744 23263 12746
rect 105 12688 110 12744
rect 166 12688 23202 12744
rect 23258 12688 23263 12744
rect 105 12686 23263 12688
rect 105 12683 171 12686
rect 23197 12683 23263 12686
rect 3244 12544 3564 12545
rect 3244 12480 3252 12544
rect 3316 12480 3332 12544
rect 3396 12480 3412 12544
rect 3476 12480 3492 12544
rect 3556 12480 3564 12544
rect 3244 12479 3564 12480
rect 6244 12544 6564 12545
rect 6244 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6412 12544
rect 6476 12480 6492 12544
rect 6556 12480 6564 12544
rect 6244 12479 6564 12480
rect 9244 12544 9564 12545
rect 9244 12480 9252 12544
rect 9316 12480 9332 12544
rect 9396 12480 9412 12544
rect 9476 12480 9492 12544
rect 9556 12480 9564 12544
rect 9244 12479 9564 12480
rect 12244 12544 12564 12545
rect 12244 12480 12252 12544
rect 12316 12480 12332 12544
rect 12396 12480 12412 12544
rect 12476 12480 12492 12544
rect 12556 12480 12564 12544
rect 12244 12479 12564 12480
rect 15244 12544 15564 12545
rect 15244 12480 15252 12544
rect 15316 12480 15332 12544
rect 15396 12480 15412 12544
rect 15476 12480 15492 12544
rect 15556 12480 15564 12544
rect 15244 12479 15564 12480
rect 18244 12544 18564 12545
rect 18244 12480 18252 12544
rect 18316 12480 18332 12544
rect 18396 12480 18412 12544
rect 18476 12480 18492 12544
rect 18556 12480 18564 12544
rect 18244 12479 18564 12480
rect 21244 12544 21564 12545
rect 21244 12480 21252 12544
rect 21316 12480 21332 12544
rect 21396 12480 21412 12544
rect 21476 12480 21492 12544
rect 21556 12480 21564 12544
rect 21244 12479 21564 12480
rect 24244 12544 24564 12545
rect 24244 12480 24252 12544
rect 24316 12480 24332 12544
rect 24396 12480 24412 12544
rect 24476 12480 24492 12544
rect 24556 12480 24564 12544
rect 24244 12479 24564 12480
rect 27244 12544 27564 12545
rect 27244 12480 27252 12544
rect 27316 12480 27332 12544
rect 27396 12480 27412 12544
rect 27476 12480 27492 12544
rect 27556 12480 27564 12544
rect 27244 12479 27564 12480
rect 1744 12000 2064 12001
rect 1744 11936 1752 12000
rect 1816 11936 1832 12000
rect 1896 11936 1912 12000
rect 1976 11936 1992 12000
rect 2056 11936 2064 12000
rect 1744 11935 2064 11936
rect 4744 12000 5064 12001
rect 4744 11936 4752 12000
rect 4816 11936 4832 12000
rect 4896 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5064 12000
rect 4744 11935 5064 11936
rect 7744 12000 8064 12001
rect 7744 11936 7752 12000
rect 7816 11936 7832 12000
rect 7896 11936 7912 12000
rect 7976 11936 7992 12000
rect 8056 11936 8064 12000
rect 7744 11935 8064 11936
rect 10744 12000 11064 12001
rect 10744 11936 10752 12000
rect 10816 11936 10832 12000
rect 10896 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11064 12000
rect 10744 11935 11064 11936
rect 13744 12000 14064 12001
rect 13744 11936 13752 12000
rect 13816 11936 13832 12000
rect 13896 11936 13912 12000
rect 13976 11936 13992 12000
rect 14056 11936 14064 12000
rect 13744 11935 14064 11936
rect 16744 12000 17064 12001
rect 16744 11936 16752 12000
rect 16816 11936 16832 12000
rect 16896 11936 16912 12000
rect 16976 11936 16992 12000
rect 17056 11936 17064 12000
rect 16744 11935 17064 11936
rect 19744 12000 20064 12001
rect 19744 11936 19752 12000
rect 19816 11936 19832 12000
rect 19896 11936 19912 12000
rect 19976 11936 19992 12000
rect 20056 11936 20064 12000
rect 19744 11935 20064 11936
rect 22744 12000 23064 12001
rect 22744 11936 22752 12000
rect 22816 11936 22832 12000
rect 22896 11936 22912 12000
rect 22976 11936 22992 12000
rect 23056 11936 23064 12000
rect 22744 11935 23064 11936
rect 25744 12000 26064 12001
rect 25744 11936 25752 12000
rect 25816 11936 25832 12000
rect 25896 11936 25912 12000
rect 25976 11936 25992 12000
rect 26056 11936 26064 12000
rect 25744 11935 26064 11936
rect 3244 11456 3564 11457
rect 3244 11392 3252 11456
rect 3316 11392 3332 11456
rect 3396 11392 3412 11456
rect 3476 11392 3492 11456
rect 3556 11392 3564 11456
rect 3244 11391 3564 11392
rect 6244 11456 6564 11457
rect 6244 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6412 11456
rect 6476 11392 6492 11456
rect 6556 11392 6564 11456
rect 6244 11391 6564 11392
rect 9244 11456 9564 11457
rect 9244 11392 9252 11456
rect 9316 11392 9332 11456
rect 9396 11392 9412 11456
rect 9476 11392 9492 11456
rect 9556 11392 9564 11456
rect 9244 11391 9564 11392
rect 12244 11456 12564 11457
rect 12244 11392 12252 11456
rect 12316 11392 12332 11456
rect 12396 11392 12412 11456
rect 12476 11392 12492 11456
rect 12556 11392 12564 11456
rect 12244 11391 12564 11392
rect 15244 11456 15564 11457
rect 15244 11392 15252 11456
rect 15316 11392 15332 11456
rect 15396 11392 15412 11456
rect 15476 11392 15492 11456
rect 15556 11392 15564 11456
rect 15244 11391 15564 11392
rect 18244 11456 18564 11457
rect 18244 11392 18252 11456
rect 18316 11392 18332 11456
rect 18396 11392 18412 11456
rect 18476 11392 18492 11456
rect 18556 11392 18564 11456
rect 18244 11391 18564 11392
rect 21244 11456 21564 11457
rect 21244 11392 21252 11456
rect 21316 11392 21332 11456
rect 21396 11392 21412 11456
rect 21476 11392 21492 11456
rect 21556 11392 21564 11456
rect 21244 11391 21564 11392
rect 24244 11456 24564 11457
rect 24244 11392 24252 11456
rect 24316 11392 24332 11456
rect 24396 11392 24412 11456
rect 24476 11392 24492 11456
rect 24556 11392 24564 11456
rect 24244 11391 24564 11392
rect 27244 11456 27564 11457
rect 27244 11392 27252 11456
rect 27316 11392 27332 11456
rect 27396 11392 27412 11456
rect 27476 11392 27492 11456
rect 27556 11392 27564 11456
rect 27244 11391 27564 11392
rect 28727 11117 29527 11144
rect 28717 11114 29527 11117
rect 28636 11112 29527 11114
rect 28636 11056 28722 11112
rect 28778 11056 29527 11112
rect 28636 11054 29527 11056
rect 28717 11051 29527 11054
rect 28727 11024 29527 11051
rect 1744 10912 2064 10913
rect 1744 10848 1752 10912
rect 1816 10848 1832 10912
rect 1896 10848 1912 10912
rect 1976 10848 1992 10912
rect 2056 10848 2064 10912
rect 1744 10847 2064 10848
rect 4744 10912 5064 10913
rect 4744 10848 4752 10912
rect 4816 10848 4832 10912
rect 4896 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5064 10912
rect 4744 10847 5064 10848
rect 7744 10912 8064 10913
rect 7744 10848 7752 10912
rect 7816 10848 7832 10912
rect 7896 10848 7912 10912
rect 7976 10848 7992 10912
rect 8056 10848 8064 10912
rect 7744 10847 8064 10848
rect 10744 10912 11064 10913
rect 10744 10848 10752 10912
rect 10816 10848 10832 10912
rect 10896 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11064 10912
rect 10744 10847 11064 10848
rect 13744 10912 14064 10913
rect 13744 10848 13752 10912
rect 13816 10848 13832 10912
rect 13896 10848 13912 10912
rect 13976 10848 13992 10912
rect 14056 10848 14064 10912
rect 13744 10847 14064 10848
rect 16744 10912 17064 10913
rect 16744 10848 16752 10912
rect 16816 10848 16832 10912
rect 16896 10848 16912 10912
rect 16976 10848 16992 10912
rect 17056 10848 17064 10912
rect 16744 10847 17064 10848
rect 19744 10912 20064 10913
rect 19744 10848 19752 10912
rect 19816 10848 19832 10912
rect 19896 10848 19912 10912
rect 19976 10848 19992 10912
rect 20056 10848 20064 10912
rect 19744 10847 20064 10848
rect 22744 10912 23064 10913
rect 22744 10848 22752 10912
rect 22816 10848 22832 10912
rect 22896 10848 22912 10912
rect 22976 10848 22992 10912
rect 23056 10848 23064 10912
rect 22744 10847 23064 10848
rect 25744 10912 26064 10913
rect 25744 10848 25752 10912
rect 25816 10848 25832 10912
rect 25896 10848 25912 10912
rect 25976 10848 25992 10912
rect 26056 10848 26064 10912
rect 25744 10847 26064 10848
rect 3244 10368 3564 10369
rect 3244 10304 3252 10368
rect 3316 10304 3332 10368
rect 3396 10304 3412 10368
rect 3476 10304 3492 10368
rect 3556 10304 3564 10368
rect 3244 10303 3564 10304
rect 6244 10368 6564 10369
rect 6244 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6412 10368
rect 6476 10304 6492 10368
rect 6556 10304 6564 10368
rect 6244 10303 6564 10304
rect 9244 10368 9564 10369
rect 9244 10304 9252 10368
rect 9316 10304 9332 10368
rect 9396 10304 9412 10368
rect 9476 10304 9492 10368
rect 9556 10304 9564 10368
rect 9244 10303 9564 10304
rect 12244 10368 12564 10369
rect 12244 10304 12252 10368
rect 12316 10304 12332 10368
rect 12396 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12564 10368
rect 12244 10303 12564 10304
rect 15244 10368 15564 10369
rect 15244 10304 15252 10368
rect 15316 10304 15332 10368
rect 15396 10304 15412 10368
rect 15476 10304 15492 10368
rect 15556 10304 15564 10368
rect 15244 10303 15564 10304
rect 18244 10368 18564 10369
rect 18244 10304 18252 10368
rect 18316 10304 18332 10368
rect 18396 10304 18412 10368
rect 18476 10304 18492 10368
rect 18556 10304 18564 10368
rect 18244 10303 18564 10304
rect 21244 10368 21564 10369
rect 21244 10304 21252 10368
rect 21316 10304 21332 10368
rect 21396 10304 21412 10368
rect 21476 10304 21492 10368
rect 21556 10304 21564 10368
rect 21244 10303 21564 10304
rect 24244 10368 24564 10369
rect 24244 10304 24252 10368
rect 24316 10304 24332 10368
rect 24396 10304 24412 10368
rect 24476 10304 24492 10368
rect 24556 10304 24564 10368
rect 24244 10303 24564 10304
rect 27244 10368 27564 10369
rect 27244 10304 27252 10368
rect 27316 10304 27332 10368
rect 27396 10304 27412 10368
rect 27476 10304 27492 10368
rect 27556 10304 27564 10368
rect 27244 10303 27564 10304
rect 19374 9964 19380 10028
rect 19444 10026 19450 10028
rect 20989 10026 21055 10029
rect 19444 10024 21055 10026
rect 19444 9968 20994 10024
rect 21050 9968 21055 10024
rect 19444 9966 21055 9968
rect 19444 9964 19450 9966
rect 20989 9963 21055 9966
rect 1744 9824 2064 9825
rect 1744 9760 1752 9824
rect 1816 9760 1832 9824
rect 1896 9760 1912 9824
rect 1976 9760 1992 9824
rect 2056 9760 2064 9824
rect 1744 9759 2064 9760
rect 4744 9824 5064 9825
rect 4744 9760 4752 9824
rect 4816 9760 4832 9824
rect 4896 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5064 9824
rect 4744 9759 5064 9760
rect 7744 9824 8064 9825
rect 7744 9760 7752 9824
rect 7816 9760 7832 9824
rect 7896 9760 7912 9824
rect 7976 9760 7992 9824
rect 8056 9760 8064 9824
rect 7744 9759 8064 9760
rect 10744 9824 11064 9825
rect 10744 9760 10752 9824
rect 10816 9760 10832 9824
rect 10896 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11064 9824
rect 10744 9759 11064 9760
rect 13744 9824 14064 9825
rect 13744 9760 13752 9824
rect 13816 9760 13832 9824
rect 13896 9760 13912 9824
rect 13976 9760 13992 9824
rect 14056 9760 14064 9824
rect 13744 9759 14064 9760
rect 16744 9824 17064 9825
rect 16744 9760 16752 9824
rect 16816 9760 16832 9824
rect 16896 9760 16912 9824
rect 16976 9760 16992 9824
rect 17056 9760 17064 9824
rect 16744 9759 17064 9760
rect 19744 9824 20064 9825
rect 19744 9760 19752 9824
rect 19816 9760 19832 9824
rect 19896 9760 19912 9824
rect 19976 9760 19992 9824
rect 20056 9760 20064 9824
rect 19744 9759 20064 9760
rect 22744 9824 23064 9825
rect 22744 9760 22752 9824
rect 22816 9760 22832 9824
rect 22896 9760 22912 9824
rect 22976 9760 22992 9824
rect 23056 9760 23064 9824
rect 22744 9759 23064 9760
rect 25744 9824 26064 9825
rect 25744 9760 25752 9824
rect 25816 9760 25832 9824
rect 25896 9760 25912 9824
rect 25976 9760 25992 9824
rect 26056 9760 26064 9824
rect 25744 9759 26064 9760
rect 3244 9280 3564 9281
rect 3244 9216 3252 9280
rect 3316 9216 3332 9280
rect 3396 9216 3412 9280
rect 3476 9216 3492 9280
rect 3556 9216 3564 9280
rect 3244 9215 3564 9216
rect 6244 9280 6564 9281
rect 6244 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6412 9280
rect 6476 9216 6492 9280
rect 6556 9216 6564 9280
rect 6244 9215 6564 9216
rect 9244 9280 9564 9281
rect 9244 9216 9252 9280
rect 9316 9216 9332 9280
rect 9396 9216 9412 9280
rect 9476 9216 9492 9280
rect 9556 9216 9564 9280
rect 9244 9215 9564 9216
rect 12244 9280 12564 9281
rect 12244 9216 12252 9280
rect 12316 9216 12332 9280
rect 12396 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12564 9280
rect 12244 9215 12564 9216
rect 15244 9280 15564 9281
rect 15244 9216 15252 9280
rect 15316 9216 15332 9280
rect 15396 9216 15412 9280
rect 15476 9216 15492 9280
rect 15556 9216 15564 9280
rect 15244 9215 15564 9216
rect 18244 9280 18564 9281
rect 18244 9216 18252 9280
rect 18316 9216 18332 9280
rect 18396 9216 18412 9280
rect 18476 9216 18492 9280
rect 18556 9216 18564 9280
rect 18244 9215 18564 9216
rect 21244 9280 21564 9281
rect 21244 9216 21252 9280
rect 21316 9216 21332 9280
rect 21396 9216 21412 9280
rect 21476 9216 21492 9280
rect 21556 9216 21564 9280
rect 21244 9215 21564 9216
rect 24244 9280 24564 9281
rect 24244 9216 24252 9280
rect 24316 9216 24332 9280
rect 24396 9216 24412 9280
rect 24476 9216 24492 9280
rect 24556 9216 24564 9280
rect 24244 9215 24564 9216
rect 27244 9280 27564 9281
rect 27244 9216 27252 9280
rect 27316 9216 27332 9280
rect 27396 9216 27412 9280
rect 27476 9216 27492 9280
rect 27556 9216 27564 9280
rect 27244 9215 27564 9216
rect 1744 8736 2064 8737
rect 1744 8672 1752 8736
rect 1816 8672 1832 8736
rect 1896 8672 1912 8736
rect 1976 8672 1992 8736
rect 2056 8672 2064 8736
rect 1744 8671 2064 8672
rect 4744 8736 5064 8737
rect 4744 8672 4752 8736
rect 4816 8672 4832 8736
rect 4896 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5064 8736
rect 4744 8671 5064 8672
rect 7744 8736 8064 8737
rect 7744 8672 7752 8736
rect 7816 8672 7832 8736
rect 7896 8672 7912 8736
rect 7976 8672 7992 8736
rect 8056 8672 8064 8736
rect 7744 8671 8064 8672
rect 10744 8736 11064 8737
rect 10744 8672 10752 8736
rect 10816 8672 10832 8736
rect 10896 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11064 8736
rect 10744 8671 11064 8672
rect 13744 8736 14064 8737
rect 13744 8672 13752 8736
rect 13816 8672 13832 8736
rect 13896 8672 13912 8736
rect 13976 8672 13992 8736
rect 14056 8672 14064 8736
rect 13744 8671 14064 8672
rect 16744 8736 17064 8737
rect 16744 8672 16752 8736
rect 16816 8672 16832 8736
rect 16896 8672 16912 8736
rect 16976 8672 16992 8736
rect 17056 8672 17064 8736
rect 16744 8671 17064 8672
rect 19744 8736 20064 8737
rect 19744 8672 19752 8736
rect 19816 8672 19832 8736
rect 19896 8672 19912 8736
rect 19976 8672 19992 8736
rect 20056 8672 20064 8736
rect 19744 8671 20064 8672
rect 22744 8736 23064 8737
rect 22744 8672 22752 8736
rect 22816 8672 22832 8736
rect 22896 8672 22912 8736
rect 22976 8672 22992 8736
rect 23056 8672 23064 8736
rect 22744 8671 23064 8672
rect 25744 8736 26064 8737
rect 25744 8672 25752 8736
rect 25816 8672 25832 8736
rect 25896 8672 25912 8736
rect 25976 8672 25992 8736
rect 26056 8672 26064 8736
rect 25744 8671 26064 8672
rect 3244 8192 3564 8193
rect 3244 8128 3252 8192
rect 3316 8128 3332 8192
rect 3396 8128 3412 8192
rect 3476 8128 3492 8192
rect 3556 8128 3564 8192
rect 3244 8127 3564 8128
rect 6244 8192 6564 8193
rect 6244 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6412 8192
rect 6476 8128 6492 8192
rect 6556 8128 6564 8192
rect 6244 8127 6564 8128
rect 9244 8192 9564 8193
rect 9244 8128 9252 8192
rect 9316 8128 9332 8192
rect 9396 8128 9412 8192
rect 9476 8128 9492 8192
rect 9556 8128 9564 8192
rect 9244 8127 9564 8128
rect 12244 8192 12564 8193
rect 12244 8128 12252 8192
rect 12316 8128 12332 8192
rect 12396 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12564 8192
rect 12244 8127 12564 8128
rect 15244 8192 15564 8193
rect 15244 8128 15252 8192
rect 15316 8128 15332 8192
rect 15396 8128 15412 8192
rect 15476 8128 15492 8192
rect 15556 8128 15564 8192
rect 15244 8127 15564 8128
rect 18244 8192 18564 8193
rect 18244 8128 18252 8192
rect 18316 8128 18332 8192
rect 18396 8128 18412 8192
rect 18476 8128 18492 8192
rect 18556 8128 18564 8192
rect 18244 8127 18564 8128
rect 21244 8192 21564 8193
rect 21244 8128 21252 8192
rect 21316 8128 21332 8192
rect 21396 8128 21412 8192
rect 21476 8128 21492 8192
rect 21556 8128 21564 8192
rect 21244 8127 21564 8128
rect 24244 8192 24564 8193
rect 24244 8128 24252 8192
rect 24316 8128 24332 8192
rect 24396 8128 24412 8192
rect 24476 8128 24492 8192
rect 24556 8128 24564 8192
rect 24244 8127 24564 8128
rect 27244 8192 27564 8193
rect 27244 8128 27252 8192
rect 27316 8128 27332 8192
rect 27396 8128 27412 8192
rect 27476 8128 27492 8192
rect 27556 8128 27564 8192
rect 27244 8127 27564 8128
rect 1744 7648 2064 7649
rect 1744 7584 1752 7648
rect 1816 7584 1832 7648
rect 1896 7584 1912 7648
rect 1976 7584 1992 7648
rect 2056 7584 2064 7648
rect 1744 7583 2064 7584
rect 4744 7648 5064 7649
rect 4744 7584 4752 7648
rect 4816 7584 4832 7648
rect 4896 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5064 7648
rect 4744 7583 5064 7584
rect 7744 7648 8064 7649
rect 7744 7584 7752 7648
rect 7816 7584 7832 7648
rect 7896 7584 7912 7648
rect 7976 7584 7992 7648
rect 8056 7584 8064 7648
rect 7744 7583 8064 7584
rect 10744 7648 11064 7649
rect 10744 7584 10752 7648
rect 10816 7584 10832 7648
rect 10896 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11064 7648
rect 10744 7583 11064 7584
rect 13744 7648 14064 7649
rect 13744 7584 13752 7648
rect 13816 7584 13832 7648
rect 13896 7584 13912 7648
rect 13976 7584 13992 7648
rect 14056 7584 14064 7648
rect 13744 7583 14064 7584
rect 16744 7648 17064 7649
rect 16744 7584 16752 7648
rect 16816 7584 16832 7648
rect 16896 7584 16912 7648
rect 16976 7584 16992 7648
rect 17056 7584 17064 7648
rect 16744 7583 17064 7584
rect 19744 7648 20064 7649
rect 19744 7584 19752 7648
rect 19816 7584 19832 7648
rect 19896 7584 19912 7648
rect 19976 7584 19992 7648
rect 20056 7584 20064 7648
rect 19744 7583 20064 7584
rect 22744 7648 23064 7649
rect 22744 7584 22752 7648
rect 22816 7584 22832 7648
rect 22896 7584 22912 7648
rect 22976 7584 22992 7648
rect 23056 7584 23064 7648
rect 22744 7583 23064 7584
rect 25744 7648 26064 7649
rect 25744 7584 25752 7648
rect 25816 7584 25832 7648
rect 25896 7584 25912 7648
rect 25976 7584 25992 7648
rect 26056 7584 26064 7648
rect 25744 7583 26064 7584
rect 3244 7104 3564 7105
rect 3244 7040 3252 7104
rect 3316 7040 3332 7104
rect 3396 7040 3412 7104
rect 3476 7040 3492 7104
rect 3556 7040 3564 7104
rect 3244 7039 3564 7040
rect 6244 7104 6564 7105
rect 6244 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6412 7104
rect 6476 7040 6492 7104
rect 6556 7040 6564 7104
rect 6244 7039 6564 7040
rect 9244 7104 9564 7105
rect 9244 7040 9252 7104
rect 9316 7040 9332 7104
rect 9396 7040 9412 7104
rect 9476 7040 9492 7104
rect 9556 7040 9564 7104
rect 9244 7039 9564 7040
rect 12244 7104 12564 7105
rect 12244 7040 12252 7104
rect 12316 7040 12332 7104
rect 12396 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12564 7104
rect 12244 7039 12564 7040
rect 15244 7104 15564 7105
rect 15244 7040 15252 7104
rect 15316 7040 15332 7104
rect 15396 7040 15412 7104
rect 15476 7040 15492 7104
rect 15556 7040 15564 7104
rect 15244 7039 15564 7040
rect 18244 7104 18564 7105
rect 18244 7040 18252 7104
rect 18316 7040 18332 7104
rect 18396 7040 18412 7104
rect 18476 7040 18492 7104
rect 18556 7040 18564 7104
rect 18244 7039 18564 7040
rect 21244 7104 21564 7105
rect 21244 7040 21252 7104
rect 21316 7040 21332 7104
rect 21396 7040 21412 7104
rect 21476 7040 21492 7104
rect 21556 7040 21564 7104
rect 21244 7039 21564 7040
rect 24244 7104 24564 7105
rect 24244 7040 24252 7104
rect 24316 7040 24332 7104
rect 24396 7040 24412 7104
rect 24476 7040 24492 7104
rect 24556 7040 24564 7104
rect 24244 7039 24564 7040
rect 27244 7104 27564 7105
rect 27244 7040 27252 7104
rect 27316 7040 27332 7104
rect 27396 7040 27412 7104
rect 27476 7040 27492 7104
rect 27556 7040 27564 7104
rect 27244 7039 27564 7040
rect 1744 6560 2064 6561
rect 1744 6496 1752 6560
rect 1816 6496 1832 6560
rect 1896 6496 1912 6560
rect 1976 6496 1992 6560
rect 2056 6496 2064 6560
rect 1744 6495 2064 6496
rect 4744 6560 5064 6561
rect 4744 6496 4752 6560
rect 4816 6496 4832 6560
rect 4896 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5064 6560
rect 4744 6495 5064 6496
rect 7744 6560 8064 6561
rect 7744 6496 7752 6560
rect 7816 6496 7832 6560
rect 7896 6496 7912 6560
rect 7976 6496 7992 6560
rect 8056 6496 8064 6560
rect 7744 6495 8064 6496
rect 10744 6560 11064 6561
rect 10744 6496 10752 6560
rect 10816 6496 10832 6560
rect 10896 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11064 6560
rect 10744 6495 11064 6496
rect 13744 6560 14064 6561
rect 13744 6496 13752 6560
rect 13816 6496 13832 6560
rect 13896 6496 13912 6560
rect 13976 6496 13992 6560
rect 14056 6496 14064 6560
rect 13744 6495 14064 6496
rect 16744 6560 17064 6561
rect 16744 6496 16752 6560
rect 16816 6496 16832 6560
rect 16896 6496 16912 6560
rect 16976 6496 16992 6560
rect 17056 6496 17064 6560
rect 16744 6495 17064 6496
rect 19744 6560 20064 6561
rect 19744 6496 19752 6560
rect 19816 6496 19832 6560
rect 19896 6496 19912 6560
rect 19976 6496 19992 6560
rect 20056 6496 20064 6560
rect 19744 6495 20064 6496
rect 22744 6560 23064 6561
rect 22744 6496 22752 6560
rect 22816 6496 22832 6560
rect 22896 6496 22912 6560
rect 22976 6496 22992 6560
rect 23056 6496 23064 6560
rect 22744 6495 23064 6496
rect 25744 6560 26064 6561
rect 25744 6496 25752 6560
rect 25816 6496 25832 6560
rect 25896 6496 25912 6560
rect 25976 6496 25992 6560
rect 26056 6496 26064 6560
rect 25744 6495 26064 6496
rect 3244 6016 3564 6017
rect 3244 5952 3252 6016
rect 3316 5952 3332 6016
rect 3396 5952 3412 6016
rect 3476 5952 3492 6016
rect 3556 5952 3564 6016
rect 3244 5951 3564 5952
rect 6244 6016 6564 6017
rect 6244 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6412 6016
rect 6476 5952 6492 6016
rect 6556 5952 6564 6016
rect 6244 5951 6564 5952
rect 9244 6016 9564 6017
rect 9244 5952 9252 6016
rect 9316 5952 9332 6016
rect 9396 5952 9412 6016
rect 9476 5952 9492 6016
rect 9556 5952 9564 6016
rect 9244 5951 9564 5952
rect 12244 6016 12564 6017
rect 12244 5952 12252 6016
rect 12316 5952 12332 6016
rect 12396 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12564 6016
rect 12244 5951 12564 5952
rect 15244 6016 15564 6017
rect 15244 5952 15252 6016
rect 15316 5952 15332 6016
rect 15396 5952 15412 6016
rect 15476 5952 15492 6016
rect 15556 5952 15564 6016
rect 15244 5951 15564 5952
rect 18244 6016 18564 6017
rect 18244 5952 18252 6016
rect 18316 5952 18332 6016
rect 18396 5952 18412 6016
rect 18476 5952 18492 6016
rect 18556 5952 18564 6016
rect 18244 5951 18564 5952
rect 21244 6016 21564 6017
rect 21244 5952 21252 6016
rect 21316 5952 21332 6016
rect 21396 5952 21412 6016
rect 21476 5952 21492 6016
rect 21556 5952 21564 6016
rect 21244 5951 21564 5952
rect 24244 6016 24564 6017
rect 24244 5952 24252 6016
rect 24316 5952 24332 6016
rect 24396 5952 24412 6016
rect 24476 5952 24492 6016
rect 24556 5952 24564 6016
rect 24244 5951 24564 5952
rect 27244 6016 27564 6017
rect 27244 5952 27252 6016
rect 27316 5952 27332 6016
rect 27396 5952 27412 6016
rect 27476 5952 27492 6016
rect 27556 5952 27564 6016
rect 27244 5951 27564 5952
rect 1744 5472 2064 5473
rect 1744 5408 1752 5472
rect 1816 5408 1832 5472
rect 1896 5408 1912 5472
rect 1976 5408 1992 5472
rect 2056 5408 2064 5472
rect 1744 5407 2064 5408
rect 4744 5472 5064 5473
rect 4744 5408 4752 5472
rect 4816 5408 4832 5472
rect 4896 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5064 5472
rect 4744 5407 5064 5408
rect 7744 5472 8064 5473
rect 7744 5408 7752 5472
rect 7816 5408 7832 5472
rect 7896 5408 7912 5472
rect 7976 5408 7992 5472
rect 8056 5408 8064 5472
rect 7744 5407 8064 5408
rect 10744 5472 11064 5473
rect 10744 5408 10752 5472
rect 10816 5408 10832 5472
rect 10896 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11064 5472
rect 10744 5407 11064 5408
rect 13744 5472 14064 5473
rect 13744 5408 13752 5472
rect 13816 5408 13832 5472
rect 13896 5408 13912 5472
rect 13976 5408 13992 5472
rect 14056 5408 14064 5472
rect 13744 5407 14064 5408
rect 16744 5472 17064 5473
rect 16744 5408 16752 5472
rect 16816 5408 16832 5472
rect 16896 5408 16912 5472
rect 16976 5408 16992 5472
rect 17056 5408 17064 5472
rect 16744 5407 17064 5408
rect 19744 5472 20064 5473
rect 19744 5408 19752 5472
rect 19816 5408 19832 5472
rect 19896 5408 19912 5472
rect 19976 5408 19992 5472
rect 20056 5408 20064 5472
rect 19744 5407 20064 5408
rect 22744 5472 23064 5473
rect 22744 5408 22752 5472
rect 22816 5408 22832 5472
rect 22896 5408 22912 5472
rect 22976 5408 22992 5472
rect 23056 5408 23064 5472
rect 22744 5407 23064 5408
rect 25744 5472 26064 5473
rect 25744 5408 25752 5472
rect 25816 5408 25832 5472
rect 25896 5408 25912 5472
rect 25976 5408 25992 5472
rect 26056 5408 26064 5472
rect 25744 5407 26064 5408
rect 3244 4928 3564 4929
rect 3244 4864 3252 4928
rect 3316 4864 3332 4928
rect 3396 4864 3412 4928
rect 3476 4864 3492 4928
rect 3556 4864 3564 4928
rect 3244 4863 3564 4864
rect 6244 4928 6564 4929
rect 6244 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6412 4928
rect 6476 4864 6492 4928
rect 6556 4864 6564 4928
rect 6244 4863 6564 4864
rect 9244 4928 9564 4929
rect 9244 4864 9252 4928
rect 9316 4864 9332 4928
rect 9396 4864 9412 4928
rect 9476 4864 9492 4928
rect 9556 4864 9564 4928
rect 9244 4863 9564 4864
rect 12244 4928 12564 4929
rect 12244 4864 12252 4928
rect 12316 4864 12332 4928
rect 12396 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12564 4928
rect 12244 4863 12564 4864
rect 15244 4928 15564 4929
rect 15244 4864 15252 4928
rect 15316 4864 15332 4928
rect 15396 4864 15412 4928
rect 15476 4864 15492 4928
rect 15556 4864 15564 4928
rect 15244 4863 15564 4864
rect 18244 4928 18564 4929
rect 18244 4864 18252 4928
rect 18316 4864 18332 4928
rect 18396 4864 18412 4928
rect 18476 4864 18492 4928
rect 18556 4864 18564 4928
rect 18244 4863 18564 4864
rect 21244 4928 21564 4929
rect 21244 4864 21252 4928
rect 21316 4864 21332 4928
rect 21396 4864 21412 4928
rect 21476 4864 21492 4928
rect 21556 4864 21564 4928
rect 21244 4863 21564 4864
rect 24244 4928 24564 4929
rect 24244 4864 24252 4928
rect 24316 4864 24332 4928
rect 24396 4864 24412 4928
rect 24476 4864 24492 4928
rect 24556 4864 24564 4928
rect 24244 4863 24564 4864
rect 27244 4928 27564 4929
rect 27244 4864 27252 4928
rect 27316 4864 27332 4928
rect 27396 4864 27412 4928
rect 27476 4864 27492 4928
rect 27556 4864 27564 4928
rect 27244 4863 27564 4864
rect 1744 4384 2064 4385
rect 1744 4320 1752 4384
rect 1816 4320 1832 4384
rect 1896 4320 1912 4384
rect 1976 4320 1992 4384
rect 2056 4320 2064 4384
rect 1744 4319 2064 4320
rect 4744 4384 5064 4385
rect 4744 4320 4752 4384
rect 4816 4320 4832 4384
rect 4896 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5064 4384
rect 4744 4319 5064 4320
rect 7744 4384 8064 4385
rect 7744 4320 7752 4384
rect 7816 4320 7832 4384
rect 7896 4320 7912 4384
rect 7976 4320 7992 4384
rect 8056 4320 8064 4384
rect 7744 4319 8064 4320
rect 10744 4384 11064 4385
rect 10744 4320 10752 4384
rect 10816 4320 10832 4384
rect 10896 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11064 4384
rect 10744 4319 11064 4320
rect 13744 4384 14064 4385
rect 13744 4320 13752 4384
rect 13816 4320 13832 4384
rect 13896 4320 13912 4384
rect 13976 4320 13992 4384
rect 14056 4320 14064 4384
rect 13744 4319 14064 4320
rect 16744 4384 17064 4385
rect 16744 4320 16752 4384
rect 16816 4320 16832 4384
rect 16896 4320 16912 4384
rect 16976 4320 16992 4384
rect 17056 4320 17064 4384
rect 16744 4319 17064 4320
rect 19744 4384 20064 4385
rect 19744 4320 19752 4384
rect 19816 4320 19832 4384
rect 19896 4320 19912 4384
rect 19976 4320 19992 4384
rect 20056 4320 20064 4384
rect 19744 4319 20064 4320
rect 22744 4384 23064 4385
rect 22744 4320 22752 4384
rect 22816 4320 22832 4384
rect 22896 4320 22912 4384
rect 22976 4320 22992 4384
rect 23056 4320 23064 4384
rect 22744 4319 23064 4320
rect 25744 4384 26064 4385
rect 25744 4320 25752 4384
rect 25816 4320 25832 4384
rect 25896 4320 25912 4384
rect 25976 4320 25992 4384
rect 26056 4320 26064 4384
rect 25744 4319 26064 4320
rect 8845 4178 8911 4181
rect 11789 4178 11855 4181
rect 12065 4178 12131 4181
rect 8845 4176 12131 4178
rect 8845 4120 8850 4176
rect 8906 4120 11794 4176
rect 11850 4120 12070 4176
rect 12126 4120 12131 4176
rect 8845 4118 12131 4120
rect 8845 4115 8911 4118
rect 11789 4115 11855 4118
rect 12065 4115 12131 4118
rect 8753 4042 8819 4045
rect 9949 4042 10015 4045
rect 8753 4040 10015 4042
rect 8753 3984 8758 4040
rect 8814 3984 9954 4040
rect 10010 3984 10015 4040
rect 8753 3982 10015 3984
rect 8753 3979 8819 3982
rect 9949 3979 10015 3982
rect 3244 3840 3564 3841
rect 3244 3776 3252 3840
rect 3316 3776 3332 3840
rect 3396 3776 3412 3840
rect 3476 3776 3492 3840
rect 3556 3776 3564 3840
rect 3244 3775 3564 3776
rect 6244 3840 6564 3841
rect 6244 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6412 3840
rect 6476 3776 6492 3840
rect 6556 3776 6564 3840
rect 6244 3775 6564 3776
rect 9244 3840 9564 3841
rect 9244 3776 9252 3840
rect 9316 3776 9332 3840
rect 9396 3776 9412 3840
rect 9476 3776 9492 3840
rect 9556 3776 9564 3840
rect 9244 3775 9564 3776
rect 12244 3840 12564 3841
rect 12244 3776 12252 3840
rect 12316 3776 12332 3840
rect 12396 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12564 3840
rect 12244 3775 12564 3776
rect 15244 3840 15564 3841
rect 15244 3776 15252 3840
rect 15316 3776 15332 3840
rect 15396 3776 15412 3840
rect 15476 3776 15492 3840
rect 15556 3776 15564 3840
rect 15244 3775 15564 3776
rect 18244 3840 18564 3841
rect 18244 3776 18252 3840
rect 18316 3776 18332 3840
rect 18396 3776 18412 3840
rect 18476 3776 18492 3840
rect 18556 3776 18564 3840
rect 18244 3775 18564 3776
rect 21244 3840 21564 3841
rect 21244 3776 21252 3840
rect 21316 3776 21332 3840
rect 21396 3776 21412 3840
rect 21476 3776 21492 3840
rect 21556 3776 21564 3840
rect 21244 3775 21564 3776
rect 24244 3840 24564 3841
rect 24244 3776 24252 3840
rect 24316 3776 24332 3840
rect 24396 3776 24412 3840
rect 24476 3776 24492 3840
rect 24556 3776 24564 3840
rect 24244 3775 24564 3776
rect 27244 3840 27564 3841
rect 27244 3776 27252 3840
rect 27316 3776 27332 3840
rect 27396 3776 27412 3840
rect 27476 3776 27492 3840
rect 27556 3776 27564 3840
rect 27244 3775 27564 3776
rect 1744 3296 2064 3297
rect 1744 3232 1752 3296
rect 1816 3232 1832 3296
rect 1896 3232 1912 3296
rect 1976 3232 1992 3296
rect 2056 3232 2064 3296
rect 1744 3231 2064 3232
rect 4744 3296 5064 3297
rect 4744 3232 4752 3296
rect 4816 3232 4832 3296
rect 4896 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5064 3296
rect 4744 3231 5064 3232
rect 7744 3296 8064 3297
rect 7744 3232 7752 3296
rect 7816 3232 7832 3296
rect 7896 3232 7912 3296
rect 7976 3232 7992 3296
rect 8056 3232 8064 3296
rect 7744 3231 8064 3232
rect 10744 3296 11064 3297
rect 10744 3232 10752 3296
rect 10816 3232 10832 3296
rect 10896 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11064 3296
rect 10744 3231 11064 3232
rect 13744 3296 14064 3297
rect 13744 3232 13752 3296
rect 13816 3232 13832 3296
rect 13896 3232 13912 3296
rect 13976 3232 13992 3296
rect 14056 3232 14064 3296
rect 13744 3231 14064 3232
rect 16744 3296 17064 3297
rect 16744 3232 16752 3296
rect 16816 3232 16832 3296
rect 16896 3232 16912 3296
rect 16976 3232 16992 3296
rect 17056 3232 17064 3296
rect 16744 3231 17064 3232
rect 19744 3296 20064 3297
rect 19744 3232 19752 3296
rect 19816 3232 19832 3296
rect 19896 3232 19912 3296
rect 19976 3232 19992 3296
rect 20056 3232 20064 3296
rect 19744 3231 20064 3232
rect 22744 3296 23064 3297
rect 22744 3232 22752 3296
rect 22816 3232 22832 3296
rect 22896 3232 22912 3296
rect 22976 3232 22992 3296
rect 23056 3232 23064 3296
rect 22744 3231 23064 3232
rect 25744 3296 26064 3297
rect 25744 3232 25752 3296
rect 25816 3232 25832 3296
rect 25896 3232 25912 3296
rect 25976 3232 25992 3296
rect 26056 3232 26064 3296
rect 25744 3231 26064 3232
rect 3244 2752 3564 2753
rect 3244 2688 3252 2752
rect 3316 2688 3332 2752
rect 3396 2688 3412 2752
rect 3476 2688 3492 2752
rect 3556 2688 3564 2752
rect 3244 2687 3564 2688
rect 6244 2752 6564 2753
rect 6244 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6412 2752
rect 6476 2688 6492 2752
rect 6556 2688 6564 2752
rect 6244 2687 6564 2688
rect 9244 2752 9564 2753
rect 9244 2688 9252 2752
rect 9316 2688 9332 2752
rect 9396 2688 9412 2752
rect 9476 2688 9492 2752
rect 9556 2688 9564 2752
rect 9244 2687 9564 2688
rect 12244 2752 12564 2753
rect 12244 2688 12252 2752
rect 12316 2688 12332 2752
rect 12396 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12564 2752
rect 12244 2687 12564 2688
rect 15244 2752 15564 2753
rect 15244 2688 15252 2752
rect 15316 2688 15332 2752
rect 15396 2688 15412 2752
rect 15476 2688 15492 2752
rect 15556 2688 15564 2752
rect 15244 2687 15564 2688
rect 18244 2752 18564 2753
rect 18244 2688 18252 2752
rect 18316 2688 18332 2752
rect 18396 2688 18412 2752
rect 18476 2688 18492 2752
rect 18556 2688 18564 2752
rect 18244 2687 18564 2688
rect 21244 2752 21564 2753
rect 21244 2688 21252 2752
rect 21316 2688 21332 2752
rect 21396 2688 21412 2752
rect 21476 2688 21492 2752
rect 21556 2688 21564 2752
rect 21244 2687 21564 2688
rect 24244 2752 24564 2753
rect 24244 2688 24252 2752
rect 24316 2688 24332 2752
rect 24396 2688 24412 2752
rect 24476 2688 24492 2752
rect 24556 2688 24564 2752
rect 24244 2687 24564 2688
rect 27244 2752 27564 2753
rect 27244 2688 27252 2752
rect 27316 2688 27332 2752
rect 27396 2688 27412 2752
rect 27476 2688 27492 2752
rect 27556 2688 27564 2752
rect 27244 2687 27564 2688
rect 1744 2208 2064 2209
rect 1744 2144 1752 2208
rect 1816 2144 1832 2208
rect 1896 2144 1912 2208
rect 1976 2144 1992 2208
rect 2056 2144 2064 2208
rect 1744 2143 2064 2144
rect 4744 2208 5064 2209
rect 4744 2144 4752 2208
rect 4816 2144 4832 2208
rect 4896 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5064 2208
rect 4744 2143 5064 2144
rect 7744 2208 8064 2209
rect 7744 2144 7752 2208
rect 7816 2144 7832 2208
rect 7896 2144 7912 2208
rect 7976 2144 7992 2208
rect 8056 2144 8064 2208
rect 7744 2143 8064 2144
rect 10744 2208 11064 2209
rect 10744 2144 10752 2208
rect 10816 2144 10832 2208
rect 10896 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11064 2208
rect 10744 2143 11064 2144
rect 13744 2208 14064 2209
rect 13744 2144 13752 2208
rect 13816 2144 13832 2208
rect 13896 2144 13912 2208
rect 13976 2144 13992 2208
rect 14056 2144 14064 2208
rect 13744 2143 14064 2144
rect 16744 2208 17064 2209
rect 16744 2144 16752 2208
rect 16816 2144 16832 2208
rect 16896 2144 16912 2208
rect 16976 2144 16992 2208
rect 17056 2144 17064 2208
rect 16744 2143 17064 2144
rect 19744 2208 20064 2209
rect 19744 2144 19752 2208
rect 19816 2144 19832 2208
rect 19896 2144 19912 2208
rect 19976 2144 19992 2208
rect 20056 2144 20064 2208
rect 19744 2143 20064 2144
rect 22744 2208 23064 2209
rect 22744 2144 22752 2208
rect 22816 2144 22832 2208
rect 22896 2144 22912 2208
rect 22976 2144 22992 2208
rect 23056 2144 23064 2208
rect 22744 2143 23064 2144
rect 25744 2208 26064 2209
rect 25744 2144 25752 2208
rect 25816 2144 25832 2208
rect 25896 2144 25912 2208
rect 25976 2144 25992 2208
rect 26056 2144 26064 2208
rect 25744 2143 26064 2144
<< via3 >>
rect 1752 29404 1816 29408
rect 1752 29348 1756 29404
rect 1756 29348 1812 29404
rect 1812 29348 1816 29404
rect 1752 29344 1816 29348
rect 1832 29404 1896 29408
rect 1832 29348 1836 29404
rect 1836 29348 1892 29404
rect 1892 29348 1896 29404
rect 1832 29344 1896 29348
rect 1912 29404 1976 29408
rect 1912 29348 1916 29404
rect 1916 29348 1972 29404
rect 1972 29348 1976 29404
rect 1912 29344 1976 29348
rect 1992 29404 2056 29408
rect 1992 29348 1996 29404
rect 1996 29348 2052 29404
rect 2052 29348 2056 29404
rect 1992 29344 2056 29348
rect 4752 29404 4816 29408
rect 4752 29348 4756 29404
rect 4756 29348 4812 29404
rect 4812 29348 4816 29404
rect 4752 29344 4816 29348
rect 4832 29404 4896 29408
rect 4832 29348 4836 29404
rect 4836 29348 4892 29404
rect 4892 29348 4896 29404
rect 4832 29344 4896 29348
rect 4912 29404 4976 29408
rect 4912 29348 4916 29404
rect 4916 29348 4972 29404
rect 4972 29348 4976 29404
rect 4912 29344 4976 29348
rect 4992 29404 5056 29408
rect 4992 29348 4996 29404
rect 4996 29348 5052 29404
rect 5052 29348 5056 29404
rect 4992 29344 5056 29348
rect 7752 29404 7816 29408
rect 7752 29348 7756 29404
rect 7756 29348 7812 29404
rect 7812 29348 7816 29404
rect 7752 29344 7816 29348
rect 7832 29404 7896 29408
rect 7832 29348 7836 29404
rect 7836 29348 7892 29404
rect 7892 29348 7896 29404
rect 7832 29344 7896 29348
rect 7912 29404 7976 29408
rect 7912 29348 7916 29404
rect 7916 29348 7972 29404
rect 7972 29348 7976 29404
rect 7912 29344 7976 29348
rect 7992 29404 8056 29408
rect 7992 29348 7996 29404
rect 7996 29348 8052 29404
rect 8052 29348 8056 29404
rect 7992 29344 8056 29348
rect 10752 29404 10816 29408
rect 10752 29348 10756 29404
rect 10756 29348 10812 29404
rect 10812 29348 10816 29404
rect 10752 29344 10816 29348
rect 10832 29404 10896 29408
rect 10832 29348 10836 29404
rect 10836 29348 10892 29404
rect 10892 29348 10896 29404
rect 10832 29344 10896 29348
rect 10912 29404 10976 29408
rect 10912 29348 10916 29404
rect 10916 29348 10972 29404
rect 10972 29348 10976 29404
rect 10912 29344 10976 29348
rect 10992 29404 11056 29408
rect 10992 29348 10996 29404
rect 10996 29348 11052 29404
rect 11052 29348 11056 29404
rect 10992 29344 11056 29348
rect 13752 29404 13816 29408
rect 13752 29348 13756 29404
rect 13756 29348 13812 29404
rect 13812 29348 13816 29404
rect 13752 29344 13816 29348
rect 13832 29404 13896 29408
rect 13832 29348 13836 29404
rect 13836 29348 13892 29404
rect 13892 29348 13896 29404
rect 13832 29344 13896 29348
rect 13912 29404 13976 29408
rect 13912 29348 13916 29404
rect 13916 29348 13972 29404
rect 13972 29348 13976 29404
rect 13912 29344 13976 29348
rect 13992 29404 14056 29408
rect 13992 29348 13996 29404
rect 13996 29348 14052 29404
rect 14052 29348 14056 29404
rect 13992 29344 14056 29348
rect 16752 29404 16816 29408
rect 16752 29348 16756 29404
rect 16756 29348 16812 29404
rect 16812 29348 16816 29404
rect 16752 29344 16816 29348
rect 16832 29404 16896 29408
rect 16832 29348 16836 29404
rect 16836 29348 16892 29404
rect 16892 29348 16896 29404
rect 16832 29344 16896 29348
rect 16912 29404 16976 29408
rect 16912 29348 16916 29404
rect 16916 29348 16972 29404
rect 16972 29348 16976 29404
rect 16912 29344 16976 29348
rect 16992 29404 17056 29408
rect 16992 29348 16996 29404
rect 16996 29348 17052 29404
rect 17052 29348 17056 29404
rect 16992 29344 17056 29348
rect 19752 29404 19816 29408
rect 19752 29348 19756 29404
rect 19756 29348 19812 29404
rect 19812 29348 19816 29404
rect 19752 29344 19816 29348
rect 19832 29404 19896 29408
rect 19832 29348 19836 29404
rect 19836 29348 19892 29404
rect 19892 29348 19896 29404
rect 19832 29344 19896 29348
rect 19912 29404 19976 29408
rect 19912 29348 19916 29404
rect 19916 29348 19972 29404
rect 19972 29348 19976 29404
rect 19912 29344 19976 29348
rect 19992 29404 20056 29408
rect 19992 29348 19996 29404
rect 19996 29348 20052 29404
rect 20052 29348 20056 29404
rect 19992 29344 20056 29348
rect 22752 29404 22816 29408
rect 22752 29348 22756 29404
rect 22756 29348 22812 29404
rect 22812 29348 22816 29404
rect 22752 29344 22816 29348
rect 22832 29404 22896 29408
rect 22832 29348 22836 29404
rect 22836 29348 22892 29404
rect 22892 29348 22896 29404
rect 22832 29344 22896 29348
rect 22912 29404 22976 29408
rect 22912 29348 22916 29404
rect 22916 29348 22972 29404
rect 22972 29348 22976 29404
rect 22912 29344 22976 29348
rect 22992 29404 23056 29408
rect 22992 29348 22996 29404
rect 22996 29348 23052 29404
rect 23052 29348 23056 29404
rect 22992 29344 23056 29348
rect 25752 29404 25816 29408
rect 25752 29348 25756 29404
rect 25756 29348 25812 29404
rect 25812 29348 25816 29404
rect 25752 29344 25816 29348
rect 25832 29404 25896 29408
rect 25832 29348 25836 29404
rect 25836 29348 25892 29404
rect 25892 29348 25896 29404
rect 25832 29344 25896 29348
rect 25912 29404 25976 29408
rect 25912 29348 25916 29404
rect 25916 29348 25972 29404
rect 25972 29348 25976 29404
rect 25912 29344 25976 29348
rect 25992 29404 26056 29408
rect 25992 29348 25996 29404
rect 25996 29348 26052 29404
rect 26052 29348 26056 29404
rect 25992 29344 26056 29348
rect 3252 28860 3316 28864
rect 3252 28804 3256 28860
rect 3256 28804 3312 28860
rect 3312 28804 3316 28860
rect 3252 28800 3316 28804
rect 3332 28860 3396 28864
rect 3332 28804 3336 28860
rect 3336 28804 3392 28860
rect 3392 28804 3396 28860
rect 3332 28800 3396 28804
rect 3412 28860 3476 28864
rect 3412 28804 3416 28860
rect 3416 28804 3472 28860
rect 3472 28804 3476 28860
rect 3412 28800 3476 28804
rect 3492 28860 3556 28864
rect 3492 28804 3496 28860
rect 3496 28804 3552 28860
rect 3552 28804 3556 28860
rect 3492 28800 3556 28804
rect 6252 28860 6316 28864
rect 6252 28804 6256 28860
rect 6256 28804 6312 28860
rect 6312 28804 6316 28860
rect 6252 28800 6316 28804
rect 6332 28860 6396 28864
rect 6332 28804 6336 28860
rect 6336 28804 6392 28860
rect 6392 28804 6396 28860
rect 6332 28800 6396 28804
rect 6412 28860 6476 28864
rect 6412 28804 6416 28860
rect 6416 28804 6472 28860
rect 6472 28804 6476 28860
rect 6412 28800 6476 28804
rect 6492 28860 6556 28864
rect 6492 28804 6496 28860
rect 6496 28804 6552 28860
rect 6552 28804 6556 28860
rect 6492 28800 6556 28804
rect 9252 28860 9316 28864
rect 9252 28804 9256 28860
rect 9256 28804 9312 28860
rect 9312 28804 9316 28860
rect 9252 28800 9316 28804
rect 9332 28860 9396 28864
rect 9332 28804 9336 28860
rect 9336 28804 9392 28860
rect 9392 28804 9396 28860
rect 9332 28800 9396 28804
rect 9412 28860 9476 28864
rect 9412 28804 9416 28860
rect 9416 28804 9472 28860
rect 9472 28804 9476 28860
rect 9412 28800 9476 28804
rect 9492 28860 9556 28864
rect 9492 28804 9496 28860
rect 9496 28804 9552 28860
rect 9552 28804 9556 28860
rect 9492 28800 9556 28804
rect 12252 28860 12316 28864
rect 12252 28804 12256 28860
rect 12256 28804 12312 28860
rect 12312 28804 12316 28860
rect 12252 28800 12316 28804
rect 12332 28860 12396 28864
rect 12332 28804 12336 28860
rect 12336 28804 12392 28860
rect 12392 28804 12396 28860
rect 12332 28800 12396 28804
rect 12412 28860 12476 28864
rect 12412 28804 12416 28860
rect 12416 28804 12472 28860
rect 12472 28804 12476 28860
rect 12412 28800 12476 28804
rect 12492 28860 12556 28864
rect 12492 28804 12496 28860
rect 12496 28804 12552 28860
rect 12552 28804 12556 28860
rect 12492 28800 12556 28804
rect 15252 28860 15316 28864
rect 15252 28804 15256 28860
rect 15256 28804 15312 28860
rect 15312 28804 15316 28860
rect 15252 28800 15316 28804
rect 15332 28860 15396 28864
rect 15332 28804 15336 28860
rect 15336 28804 15392 28860
rect 15392 28804 15396 28860
rect 15332 28800 15396 28804
rect 15412 28860 15476 28864
rect 15412 28804 15416 28860
rect 15416 28804 15472 28860
rect 15472 28804 15476 28860
rect 15412 28800 15476 28804
rect 15492 28860 15556 28864
rect 15492 28804 15496 28860
rect 15496 28804 15552 28860
rect 15552 28804 15556 28860
rect 15492 28800 15556 28804
rect 18252 28860 18316 28864
rect 18252 28804 18256 28860
rect 18256 28804 18312 28860
rect 18312 28804 18316 28860
rect 18252 28800 18316 28804
rect 18332 28860 18396 28864
rect 18332 28804 18336 28860
rect 18336 28804 18392 28860
rect 18392 28804 18396 28860
rect 18332 28800 18396 28804
rect 18412 28860 18476 28864
rect 18412 28804 18416 28860
rect 18416 28804 18472 28860
rect 18472 28804 18476 28860
rect 18412 28800 18476 28804
rect 18492 28860 18556 28864
rect 18492 28804 18496 28860
rect 18496 28804 18552 28860
rect 18552 28804 18556 28860
rect 18492 28800 18556 28804
rect 21252 28860 21316 28864
rect 21252 28804 21256 28860
rect 21256 28804 21312 28860
rect 21312 28804 21316 28860
rect 21252 28800 21316 28804
rect 21332 28860 21396 28864
rect 21332 28804 21336 28860
rect 21336 28804 21392 28860
rect 21392 28804 21396 28860
rect 21332 28800 21396 28804
rect 21412 28860 21476 28864
rect 21412 28804 21416 28860
rect 21416 28804 21472 28860
rect 21472 28804 21476 28860
rect 21412 28800 21476 28804
rect 21492 28860 21556 28864
rect 21492 28804 21496 28860
rect 21496 28804 21552 28860
rect 21552 28804 21556 28860
rect 21492 28800 21556 28804
rect 24252 28860 24316 28864
rect 24252 28804 24256 28860
rect 24256 28804 24312 28860
rect 24312 28804 24316 28860
rect 24252 28800 24316 28804
rect 24332 28860 24396 28864
rect 24332 28804 24336 28860
rect 24336 28804 24392 28860
rect 24392 28804 24396 28860
rect 24332 28800 24396 28804
rect 24412 28860 24476 28864
rect 24412 28804 24416 28860
rect 24416 28804 24472 28860
rect 24472 28804 24476 28860
rect 24412 28800 24476 28804
rect 24492 28860 24556 28864
rect 24492 28804 24496 28860
rect 24496 28804 24552 28860
rect 24552 28804 24556 28860
rect 24492 28800 24556 28804
rect 27252 28860 27316 28864
rect 27252 28804 27256 28860
rect 27256 28804 27312 28860
rect 27312 28804 27316 28860
rect 27252 28800 27316 28804
rect 27332 28860 27396 28864
rect 27332 28804 27336 28860
rect 27336 28804 27392 28860
rect 27392 28804 27396 28860
rect 27332 28800 27396 28804
rect 27412 28860 27476 28864
rect 27412 28804 27416 28860
rect 27416 28804 27472 28860
rect 27472 28804 27476 28860
rect 27412 28800 27476 28804
rect 27492 28860 27556 28864
rect 27492 28804 27496 28860
rect 27496 28804 27552 28860
rect 27552 28804 27556 28860
rect 27492 28800 27556 28804
rect 1752 28316 1816 28320
rect 1752 28260 1756 28316
rect 1756 28260 1812 28316
rect 1812 28260 1816 28316
rect 1752 28256 1816 28260
rect 1832 28316 1896 28320
rect 1832 28260 1836 28316
rect 1836 28260 1892 28316
rect 1892 28260 1896 28316
rect 1832 28256 1896 28260
rect 1912 28316 1976 28320
rect 1912 28260 1916 28316
rect 1916 28260 1972 28316
rect 1972 28260 1976 28316
rect 1912 28256 1976 28260
rect 1992 28316 2056 28320
rect 1992 28260 1996 28316
rect 1996 28260 2052 28316
rect 2052 28260 2056 28316
rect 1992 28256 2056 28260
rect 4752 28316 4816 28320
rect 4752 28260 4756 28316
rect 4756 28260 4812 28316
rect 4812 28260 4816 28316
rect 4752 28256 4816 28260
rect 4832 28316 4896 28320
rect 4832 28260 4836 28316
rect 4836 28260 4892 28316
rect 4892 28260 4896 28316
rect 4832 28256 4896 28260
rect 4912 28316 4976 28320
rect 4912 28260 4916 28316
rect 4916 28260 4972 28316
rect 4972 28260 4976 28316
rect 4912 28256 4976 28260
rect 4992 28316 5056 28320
rect 4992 28260 4996 28316
rect 4996 28260 5052 28316
rect 5052 28260 5056 28316
rect 4992 28256 5056 28260
rect 7752 28316 7816 28320
rect 7752 28260 7756 28316
rect 7756 28260 7812 28316
rect 7812 28260 7816 28316
rect 7752 28256 7816 28260
rect 7832 28316 7896 28320
rect 7832 28260 7836 28316
rect 7836 28260 7892 28316
rect 7892 28260 7896 28316
rect 7832 28256 7896 28260
rect 7912 28316 7976 28320
rect 7912 28260 7916 28316
rect 7916 28260 7972 28316
rect 7972 28260 7976 28316
rect 7912 28256 7976 28260
rect 7992 28316 8056 28320
rect 7992 28260 7996 28316
rect 7996 28260 8052 28316
rect 8052 28260 8056 28316
rect 7992 28256 8056 28260
rect 10752 28316 10816 28320
rect 10752 28260 10756 28316
rect 10756 28260 10812 28316
rect 10812 28260 10816 28316
rect 10752 28256 10816 28260
rect 10832 28316 10896 28320
rect 10832 28260 10836 28316
rect 10836 28260 10892 28316
rect 10892 28260 10896 28316
rect 10832 28256 10896 28260
rect 10912 28316 10976 28320
rect 10912 28260 10916 28316
rect 10916 28260 10972 28316
rect 10972 28260 10976 28316
rect 10912 28256 10976 28260
rect 10992 28316 11056 28320
rect 10992 28260 10996 28316
rect 10996 28260 11052 28316
rect 11052 28260 11056 28316
rect 10992 28256 11056 28260
rect 13752 28316 13816 28320
rect 13752 28260 13756 28316
rect 13756 28260 13812 28316
rect 13812 28260 13816 28316
rect 13752 28256 13816 28260
rect 13832 28316 13896 28320
rect 13832 28260 13836 28316
rect 13836 28260 13892 28316
rect 13892 28260 13896 28316
rect 13832 28256 13896 28260
rect 13912 28316 13976 28320
rect 13912 28260 13916 28316
rect 13916 28260 13972 28316
rect 13972 28260 13976 28316
rect 13912 28256 13976 28260
rect 13992 28316 14056 28320
rect 13992 28260 13996 28316
rect 13996 28260 14052 28316
rect 14052 28260 14056 28316
rect 13992 28256 14056 28260
rect 16752 28316 16816 28320
rect 16752 28260 16756 28316
rect 16756 28260 16812 28316
rect 16812 28260 16816 28316
rect 16752 28256 16816 28260
rect 16832 28316 16896 28320
rect 16832 28260 16836 28316
rect 16836 28260 16892 28316
rect 16892 28260 16896 28316
rect 16832 28256 16896 28260
rect 16912 28316 16976 28320
rect 16912 28260 16916 28316
rect 16916 28260 16972 28316
rect 16972 28260 16976 28316
rect 16912 28256 16976 28260
rect 16992 28316 17056 28320
rect 16992 28260 16996 28316
rect 16996 28260 17052 28316
rect 17052 28260 17056 28316
rect 16992 28256 17056 28260
rect 19752 28316 19816 28320
rect 19752 28260 19756 28316
rect 19756 28260 19812 28316
rect 19812 28260 19816 28316
rect 19752 28256 19816 28260
rect 19832 28316 19896 28320
rect 19832 28260 19836 28316
rect 19836 28260 19892 28316
rect 19892 28260 19896 28316
rect 19832 28256 19896 28260
rect 19912 28316 19976 28320
rect 19912 28260 19916 28316
rect 19916 28260 19972 28316
rect 19972 28260 19976 28316
rect 19912 28256 19976 28260
rect 19992 28316 20056 28320
rect 19992 28260 19996 28316
rect 19996 28260 20052 28316
rect 20052 28260 20056 28316
rect 19992 28256 20056 28260
rect 22752 28316 22816 28320
rect 22752 28260 22756 28316
rect 22756 28260 22812 28316
rect 22812 28260 22816 28316
rect 22752 28256 22816 28260
rect 22832 28316 22896 28320
rect 22832 28260 22836 28316
rect 22836 28260 22892 28316
rect 22892 28260 22896 28316
rect 22832 28256 22896 28260
rect 22912 28316 22976 28320
rect 22912 28260 22916 28316
rect 22916 28260 22972 28316
rect 22972 28260 22976 28316
rect 22912 28256 22976 28260
rect 22992 28316 23056 28320
rect 22992 28260 22996 28316
rect 22996 28260 23052 28316
rect 23052 28260 23056 28316
rect 22992 28256 23056 28260
rect 25752 28316 25816 28320
rect 25752 28260 25756 28316
rect 25756 28260 25812 28316
rect 25812 28260 25816 28316
rect 25752 28256 25816 28260
rect 25832 28316 25896 28320
rect 25832 28260 25836 28316
rect 25836 28260 25892 28316
rect 25892 28260 25896 28316
rect 25832 28256 25896 28260
rect 25912 28316 25976 28320
rect 25912 28260 25916 28316
rect 25916 28260 25972 28316
rect 25972 28260 25976 28316
rect 25912 28256 25976 28260
rect 25992 28316 26056 28320
rect 25992 28260 25996 28316
rect 25996 28260 26052 28316
rect 26052 28260 26056 28316
rect 25992 28256 26056 28260
rect 3252 27772 3316 27776
rect 3252 27716 3256 27772
rect 3256 27716 3312 27772
rect 3312 27716 3316 27772
rect 3252 27712 3316 27716
rect 3332 27772 3396 27776
rect 3332 27716 3336 27772
rect 3336 27716 3392 27772
rect 3392 27716 3396 27772
rect 3332 27712 3396 27716
rect 3412 27772 3476 27776
rect 3412 27716 3416 27772
rect 3416 27716 3472 27772
rect 3472 27716 3476 27772
rect 3412 27712 3476 27716
rect 3492 27772 3556 27776
rect 3492 27716 3496 27772
rect 3496 27716 3552 27772
rect 3552 27716 3556 27772
rect 3492 27712 3556 27716
rect 6252 27772 6316 27776
rect 6252 27716 6256 27772
rect 6256 27716 6312 27772
rect 6312 27716 6316 27772
rect 6252 27712 6316 27716
rect 6332 27772 6396 27776
rect 6332 27716 6336 27772
rect 6336 27716 6392 27772
rect 6392 27716 6396 27772
rect 6332 27712 6396 27716
rect 6412 27772 6476 27776
rect 6412 27716 6416 27772
rect 6416 27716 6472 27772
rect 6472 27716 6476 27772
rect 6412 27712 6476 27716
rect 6492 27772 6556 27776
rect 6492 27716 6496 27772
rect 6496 27716 6552 27772
rect 6552 27716 6556 27772
rect 6492 27712 6556 27716
rect 9252 27772 9316 27776
rect 9252 27716 9256 27772
rect 9256 27716 9312 27772
rect 9312 27716 9316 27772
rect 9252 27712 9316 27716
rect 9332 27772 9396 27776
rect 9332 27716 9336 27772
rect 9336 27716 9392 27772
rect 9392 27716 9396 27772
rect 9332 27712 9396 27716
rect 9412 27772 9476 27776
rect 9412 27716 9416 27772
rect 9416 27716 9472 27772
rect 9472 27716 9476 27772
rect 9412 27712 9476 27716
rect 9492 27772 9556 27776
rect 9492 27716 9496 27772
rect 9496 27716 9552 27772
rect 9552 27716 9556 27772
rect 9492 27712 9556 27716
rect 12252 27772 12316 27776
rect 12252 27716 12256 27772
rect 12256 27716 12312 27772
rect 12312 27716 12316 27772
rect 12252 27712 12316 27716
rect 12332 27772 12396 27776
rect 12332 27716 12336 27772
rect 12336 27716 12392 27772
rect 12392 27716 12396 27772
rect 12332 27712 12396 27716
rect 12412 27772 12476 27776
rect 12412 27716 12416 27772
rect 12416 27716 12472 27772
rect 12472 27716 12476 27772
rect 12412 27712 12476 27716
rect 12492 27772 12556 27776
rect 12492 27716 12496 27772
rect 12496 27716 12552 27772
rect 12552 27716 12556 27772
rect 12492 27712 12556 27716
rect 15252 27772 15316 27776
rect 15252 27716 15256 27772
rect 15256 27716 15312 27772
rect 15312 27716 15316 27772
rect 15252 27712 15316 27716
rect 15332 27772 15396 27776
rect 15332 27716 15336 27772
rect 15336 27716 15392 27772
rect 15392 27716 15396 27772
rect 15332 27712 15396 27716
rect 15412 27772 15476 27776
rect 15412 27716 15416 27772
rect 15416 27716 15472 27772
rect 15472 27716 15476 27772
rect 15412 27712 15476 27716
rect 15492 27772 15556 27776
rect 15492 27716 15496 27772
rect 15496 27716 15552 27772
rect 15552 27716 15556 27772
rect 15492 27712 15556 27716
rect 18252 27772 18316 27776
rect 18252 27716 18256 27772
rect 18256 27716 18312 27772
rect 18312 27716 18316 27772
rect 18252 27712 18316 27716
rect 18332 27772 18396 27776
rect 18332 27716 18336 27772
rect 18336 27716 18392 27772
rect 18392 27716 18396 27772
rect 18332 27712 18396 27716
rect 18412 27772 18476 27776
rect 18412 27716 18416 27772
rect 18416 27716 18472 27772
rect 18472 27716 18476 27772
rect 18412 27712 18476 27716
rect 18492 27772 18556 27776
rect 18492 27716 18496 27772
rect 18496 27716 18552 27772
rect 18552 27716 18556 27772
rect 18492 27712 18556 27716
rect 21252 27772 21316 27776
rect 21252 27716 21256 27772
rect 21256 27716 21312 27772
rect 21312 27716 21316 27772
rect 21252 27712 21316 27716
rect 21332 27772 21396 27776
rect 21332 27716 21336 27772
rect 21336 27716 21392 27772
rect 21392 27716 21396 27772
rect 21332 27712 21396 27716
rect 21412 27772 21476 27776
rect 21412 27716 21416 27772
rect 21416 27716 21472 27772
rect 21472 27716 21476 27772
rect 21412 27712 21476 27716
rect 21492 27772 21556 27776
rect 21492 27716 21496 27772
rect 21496 27716 21552 27772
rect 21552 27716 21556 27772
rect 21492 27712 21556 27716
rect 24252 27772 24316 27776
rect 24252 27716 24256 27772
rect 24256 27716 24312 27772
rect 24312 27716 24316 27772
rect 24252 27712 24316 27716
rect 24332 27772 24396 27776
rect 24332 27716 24336 27772
rect 24336 27716 24392 27772
rect 24392 27716 24396 27772
rect 24332 27712 24396 27716
rect 24412 27772 24476 27776
rect 24412 27716 24416 27772
rect 24416 27716 24472 27772
rect 24472 27716 24476 27772
rect 24412 27712 24476 27716
rect 24492 27772 24556 27776
rect 24492 27716 24496 27772
rect 24496 27716 24552 27772
rect 24552 27716 24556 27772
rect 24492 27712 24556 27716
rect 27252 27772 27316 27776
rect 27252 27716 27256 27772
rect 27256 27716 27312 27772
rect 27312 27716 27316 27772
rect 27252 27712 27316 27716
rect 27332 27772 27396 27776
rect 27332 27716 27336 27772
rect 27336 27716 27392 27772
rect 27392 27716 27396 27772
rect 27332 27712 27396 27716
rect 27412 27772 27476 27776
rect 27412 27716 27416 27772
rect 27416 27716 27472 27772
rect 27472 27716 27476 27772
rect 27412 27712 27476 27716
rect 27492 27772 27556 27776
rect 27492 27716 27496 27772
rect 27496 27716 27552 27772
rect 27552 27716 27556 27772
rect 27492 27712 27556 27716
rect 1752 27228 1816 27232
rect 1752 27172 1756 27228
rect 1756 27172 1812 27228
rect 1812 27172 1816 27228
rect 1752 27168 1816 27172
rect 1832 27228 1896 27232
rect 1832 27172 1836 27228
rect 1836 27172 1892 27228
rect 1892 27172 1896 27228
rect 1832 27168 1896 27172
rect 1912 27228 1976 27232
rect 1912 27172 1916 27228
rect 1916 27172 1972 27228
rect 1972 27172 1976 27228
rect 1912 27168 1976 27172
rect 1992 27228 2056 27232
rect 1992 27172 1996 27228
rect 1996 27172 2052 27228
rect 2052 27172 2056 27228
rect 1992 27168 2056 27172
rect 4752 27228 4816 27232
rect 4752 27172 4756 27228
rect 4756 27172 4812 27228
rect 4812 27172 4816 27228
rect 4752 27168 4816 27172
rect 4832 27228 4896 27232
rect 4832 27172 4836 27228
rect 4836 27172 4892 27228
rect 4892 27172 4896 27228
rect 4832 27168 4896 27172
rect 4912 27228 4976 27232
rect 4912 27172 4916 27228
rect 4916 27172 4972 27228
rect 4972 27172 4976 27228
rect 4912 27168 4976 27172
rect 4992 27228 5056 27232
rect 4992 27172 4996 27228
rect 4996 27172 5052 27228
rect 5052 27172 5056 27228
rect 4992 27168 5056 27172
rect 7752 27228 7816 27232
rect 7752 27172 7756 27228
rect 7756 27172 7812 27228
rect 7812 27172 7816 27228
rect 7752 27168 7816 27172
rect 7832 27228 7896 27232
rect 7832 27172 7836 27228
rect 7836 27172 7892 27228
rect 7892 27172 7896 27228
rect 7832 27168 7896 27172
rect 7912 27228 7976 27232
rect 7912 27172 7916 27228
rect 7916 27172 7972 27228
rect 7972 27172 7976 27228
rect 7912 27168 7976 27172
rect 7992 27228 8056 27232
rect 7992 27172 7996 27228
rect 7996 27172 8052 27228
rect 8052 27172 8056 27228
rect 7992 27168 8056 27172
rect 10752 27228 10816 27232
rect 10752 27172 10756 27228
rect 10756 27172 10812 27228
rect 10812 27172 10816 27228
rect 10752 27168 10816 27172
rect 10832 27228 10896 27232
rect 10832 27172 10836 27228
rect 10836 27172 10892 27228
rect 10892 27172 10896 27228
rect 10832 27168 10896 27172
rect 10912 27228 10976 27232
rect 10912 27172 10916 27228
rect 10916 27172 10972 27228
rect 10972 27172 10976 27228
rect 10912 27168 10976 27172
rect 10992 27228 11056 27232
rect 10992 27172 10996 27228
rect 10996 27172 11052 27228
rect 11052 27172 11056 27228
rect 10992 27168 11056 27172
rect 13752 27228 13816 27232
rect 13752 27172 13756 27228
rect 13756 27172 13812 27228
rect 13812 27172 13816 27228
rect 13752 27168 13816 27172
rect 13832 27228 13896 27232
rect 13832 27172 13836 27228
rect 13836 27172 13892 27228
rect 13892 27172 13896 27228
rect 13832 27168 13896 27172
rect 13912 27228 13976 27232
rect 13912 27172 13916 27228
rect 13916 27172 13972 27228
rect 13972 27172 13976 27228
rect 13912 27168 13976 27172
rect 13992 27228 14056 27232
rect 13992 27172 13996 27228
rect 13996 27172 14052 27228
rect 14052 27172 14056 27228
rect 13992 27168 14056 27172
rect 16752 27228 16816 27232
rect 16752 27172 16756 27228
rect 16756 27172 16812 27228
rect 16812 27172 16816 27228
rect 16752 27168 16816 27172
rect 16832 27228 16896 27232
rect 16832 27172 16836 27228
rect 16836 27172 16892 27228
rect 16892 27172 16896 27228
rect 16832 27168 16896 27172
rect 16912 27228 16976 27232
rect 16912 27172 16916 27228
rect 16916 27172 16972 27228
rect 16972 27172 16976 27228
rect 16912 27168 16976 27172
rect 16992 27228 17056 27232
rect 16992 27172 16996 27228
rect 16996 27172 17052 27228
rect 17052 27172 17056 27228
rect 16992 27168 17056 27172
rect 19752 27228 19816 27232
rect 19752 27172 19756 27228
rect 19756 27172 19812 27228
rect 19812 27172 19816 27228
rect 19752 27168 19816 27172
rect 19832 27228 19896 27232
rect 19832 27172 19836 27228
rect 19836 27172 19892 27228
rect 19892 27172 19896 27228
rect 19832 27168 19896 27172
rect 19912 27228 19976 27232
rect 19912 27172 19916 27228
rect 19916 27172 19972 27228
rect 19972 27172 19976 27228
rect 19912 27168 19976 27172
rect 19992 27228 20056 27232
rect 19992 27172 19996 27228
rect 19996 27172 20052 27228
rect 20052 27172 20056 27228
rect 19992 27168 20056 27172
rect 22752 27228 22816 27232
rect 22752 27172 22756 27228
rect 22756 27172 22812 27228
rect 22812 27172 22816 27228
rect 22752 27168 22816 27172
rect 22832 27228 22896 27232
rect 22832 27172 22836 27228
rect 22836 27172 22892 27228
rect 22892 27172 22896 27228
rect 22832 27168 22896 27172
rect 22912 27228 22976 27232
rect 22912 27172 22916 27228
rect 22916 27172 22972 27228
rect 22972 27172 22976 27228
rect 22912 27168 22976 27172
rect 22992 27228 23056 27232
rect 22992 27172 22996 27228
rect 22996 27172 23052 27228
rect 23052 27172 23056 27228
rect 22992 27168 23056 27172
rect 25752 27228 25816 27232
rect 25752 27172 25756 27228
rect 25756 27172 25812 27228
rect 25812 27172 25816 27228
rect 25752 27168 25816 27172
rect 25832 27228 25896 27232
rect 25832 27172 25836 27228
rect 25836 27172 25892 27228
rect 25892 27172 25896 27228
rect 25832 27168 25896 27172
rect 25912 27228 25976 27232
rect 25912 27172 25916 27228
rect 25916 27172 25972 27228
rect 25972 27172 25976 27228
rect 25912 27168 25976 27172
rect 25992 27228 26056 27232
rect 25992 27172 25996 27228
rect 25996 27172 26052 27228
rect 26052 27172 26056 27228
rect 25992 27168 26056 27172
rect 3252 26684 3316 26688
rect 3252 26628 3256 26684
rect 3256 26628 3312 26684
rect 3312 26628 3316 26684
rect 3252 26624 3316 26628
rect 3332 26684 3396 26688
rect 3332 26628 3336 26684
rect 3336 26628 3392 26684
rect 3392 26628 3396 26684
rect 3332 26624 3396 26628
rect 3412 26684 3476 26688
rect 3412 26628 3416 26684
rect 3416 26628 3472 26684
rect 3472 26628 3476 26684
rect 3412 26624 3476 26628
rect 3492 26684 3556 26688
rect 3492 26628 3496 26684
rect 3496 26628 3552 26684
rect 3552 26628 3556 26684
rect 3492 26624 3556 26628
rect 6252 26684 6316 26688
rect 6252 26628 6256 26684
rect 6256 26628 6312 26684
rect 6312 26628 6316 26684
rect 6252 26624 6316 26628
rect 6332 26684 6396 26688
rect 6332 26628 6336 26684
rect 6336 26628 6392 26684
rect 6392 26628 6396 26684
rect 6332 26624 6396 26628
rect 6412 26684 6476 26688
rect 6412 26628 6416 26684
rect 6416 26628 6472 26684
rect 6472 26628 6476 26684
rect 6412 26624 6476 26628
rect 6492 26684 6556 26688
rect 6492 26628 6496 26684
rect 6496 26628 6552 26684
rect 6552 26628 6556 26684
rect 6492 26624 6556 26628
rect 9252 26684 9316 26688
rect 9252 26628 9256 26684
rect 9256 26628 9312 26684
rect 9312 26628 9316 26684
rect 9252 26624 9316 26628
rect 9332 26684 9396 26688
rect 9332 26628 9336 26684
rect 9336 26628 9392 26684
rect 9392 26628 9396 26684
rect 9332 26624 9396 26628
rect 9412 26684 9476 26688
rect 9412 26628 9416 26684
rect 9416 26628 9472 26684
rect 9472 26628 9476 26684
rect 9412 26624 9476 26628
rect 9492 26684 9556 26688
rect 9492 26628 9496 26684
rect 9496 26628 9552 26684
rect 9552 26628 9556 26684
rect 9492 26624 9556 26628
rect 12252 26684 12316 26688
rect 12252 26628 12256 26684
rect 12256 26628 12312 26684
rect 12312 26628 12316 26684
rect 12252 26624 12316 26628
rect 12332 26684 12396 26688
rect 12332 26628 12336 26684
rect 12336 26628 12392 26684
rect 12392 26628 12396 26684
rect 12332 26624 12396 26628
rect 12412 26684 12476 26688
rect 12412 26628 12416 26684
rect 12416 26628 12472 26684
rect 12472 26628 12476 26684
rect 12412 26624 12476 26628
rect 12492 26684 12556 26688
rect 12492 26628 12496 26684
rect 12496 26628 12552 26684
rect 12552 26628 12556 26684
rect 12492 26624 12556 26628
rect 15252 26684 15316 26688
rect 15252 26628 15256 26684
rect 15256 26628 15312 26684
rect 15312 26628 15316 26684
rect 15252 26624 15316 26628
rect 15332 26684 15396 26688
rect 15332 26628 15336 26684
rect 15336 26628 15392 26684
rect 15392 26628 15396 26684
rect 15332 26624 15396 26628
rect 15412 26684 15476 26688
rect 15412 26628 15416 26684
rect 15416 26628 15472 26684
rect 15472 26628 15476 26684
rect 15412 26624 15476 26628
rect 15492 26684 15556 26688
rect 15492 26628 15496 26684
rect 15496 26628 15552 26684
rect 15552 26628 15556 26684
rect 15492 26624 15556 26628
rect 18252 26684 18316 26688
rect 18252 26628 18256 26684
rect 18256 26628 18312 26684
rect 18312 26628 18316 26684
rect 18252 26624 18316 26628
rect 18332 26684 18396 26688
rect 18332 26628 18336 26684
rect 18336 26628 18392 26684
rect 18392 26628 18396 26684
rect 18332 26624 18396 26628
rect 18412 26684 18476 26688
rect 18412 26628 18416 26684
rect 18416 26628 18472 26684
rect 18472 26628 18476 26684
rect 18412 26624 18476 26628
rect 18492 26684 18556 26688
rect 18492 26628 18496 26684
rect 18496 26628 18552 26684
rect 18552 26628 18556 26684
rect 18492 26624 18556 26628
rect 21252 26684 21316 26688
rect 21252 26628 21256 26684
rect 21256 26628 21312 26684
rect 21312 26628 21316 26684
rect 21252 26624 21316 26628
rect 21332 26684 21396 26688
rect 21332 26628 21336 26684
rect 21336 26628 21392 26684
rect 21392 26628 21396 26684
rect 21332 26624 21396 26628
rect 21412 26684 21476 26688
rect 21412 26628 21416 26684
rect 21416 26628 21472 26684
rect 21472 26628 21476 26684
rect 21412 26624 21476 26628
rect 21492 26684 21556 26688
rect 21492 26628 21496 26684
rect 21496 26628 21552 26684
rect 21552 26628 21556 26684
rect 21492 26624 21556 26628
rect 24252 26684 24316 26688
rect 24252 26628 24256 26684
rect 24256 26628 24312 26684
rect 24312 26628 24316 26684
rect 24252 26624 24316 26628
rect 24332 26684 24396 26688
rect 24332 26628 24336 26684
rect 24336 26628 24392 26684
rect 24392 26628 24396 26684
rect 24332 26624 24396 26628
rect 24412 26684 24476 26688
rect 24412 26628 24416 26684
rect 24416 26628 24472 26684
rect 24472 26628 24476 26684
rect 24412 26624 24476 26628
rect 24492 26684 24556 26688
rect 24492 26628 24496 26684
rect 24496 26628 24552 26684
rect 24552 26628 24556 26684
rect 24492 26624 24556 26628
rect 27252 26684 27316 26688
rect 27252 26628 27256 26684
rect 27256 26628 27312 26684
rect 27312 26628 27316 26684
rect 27252 26624 27316 26628
rect 27332 26684 27396 26688
rect 27332 26628 27336 26684
rect 27336 26628 27392 26684
rect 27392 26628 27396 26684
rect 27332 26624 27396 26628
rect 27412 26684 27476 26688
rect 27412 26628 27416 26684
rect 27416 26628 27472 26684
rect 27472 26628 27476 26684
rect 27412 26624 27476 26628
rect 27492 26684 27556 26688
rect 27492 26628 27496 26684
rect 27496 26628 27552 26684
rect 27552 26628 27556 26684
rect 27492 26624 27556 26628
rect 1752 26140 1816 26144
rect 1752 26084 1756 26140
rect 1756 26084 1812 26140
rect 1812 26084 1816 26140
rect 1752 26080 1816 26084
rect 1832 26140 1896 26144
rect 1832 26084 1836 26140
rect 1836 26084 1892 26140
rect 1892 26084 1896 26140
rect 1832 26080 1896 26084
rect 1912 26140 1976 26144
rect 1912 26084 1916 26140
rect 1916 26084 1972 26140
rect 1972 26084 1976 26140
rect 1912 26080 1976 26084
rect 1992 26140 2056 26144
rect 1992 26084 1996 26140
rect 1996 26084 2052 26140
rect 2052 26084 2056 26140
rect 1992 26080 2056 26084
rect 4752 26140 4816 26144
rect 4752 26084 4756 26140
rect 4756 26084 4812 26140
rect 4812 26084 4816 26140
rect 4752 26080 4816 26084
rect 4832 26140 4896 26144
rect 4832 26084 4836 26140
rect 4836 26084 4892 26140
rect 4892 26084 4896 26140
rect 4832 26080 4896 26084
rect 4912 26140 4976 26144
rect 4912 26084 4916 26140
rect 4916 26084 4972 26140
rect 4972 26084 4976 26140
rect 4912 26080 4976 26084
rect 4992 26140 5056 26144
rect 4992 26084 4996 26140
rect 4996 26084 5052 26140
rect 5052 26084 5056 26140
rect 4992 26080 5056 26084
rect 7752 26140 7816 26144
rect 7752 26084 7756 26140
rect 7756 26084 7812 26140
rect 7812 26084 7816 26140
rect 7752 26080 7816 26084
rect 7832 26140 7896 26144
rect 7832 26084 7836 26140
rect 7836 26084 7892 26140
rect 7892 26084 7896 26140
rect 7832 26080 7896 26084
rect 7912 26140 7976 26144
rect 7912 26084 7916 26140
rect 7916 26084 7972 26140
rect 7972 26084 7976 26140
rect 7912 26080 7976 26084
rect 7992 26140 8056 26144
rect 7992 26084 7996 26140
rect 7996 26084 8052 26140
rect 8052 26084 8056 26140
rect 7992 26080 8056 26084
rect 10752 26140 10816 26144
rect 10752 26084 10756 26140
rect 10756 26084 10812 26140
rect 10812 26084 10816 26140
rect 10752 26080 10816 26084
rect 10832 26140 10896 26144
rect 10832 26084 10836 26140
rect 10836 26084 10892 26140
rect 10892 26084 10896 26140
rect 10832 26080 10896 26084
rect 10912 26140 10976 26144
rect 10912 26084 10916 26140
rect 10916 26084 10972 26140
rect 10972 26084 10976 26140
rect 10912 26080 10976 26084
rect 10992 26140 11056 26144
rect 10992 26084 10996 26140
rect 10996 26084 11052 26140
rect 11052 26084 11056 26140
rect 10992 26080 11056 26084
rect 13752 26140 13816 26144
rect 13752 26084 13756 26140
rect 13756 26084 13812 26140
rect 13812 26084 13816 26140
rect 13752 26080 13816 26084
rect 13832 26140 13896 26144
rect 13832 26084 13836 26140
rect 13836 26084 13892 26140
rect 13892 26084 13896 26140
rect 13832 26080 13896 26084
rect 13912 26140 13976 26144
rect 13912 26084 13916 26140
rect 13916 26084 13972 26140
rect 13972 26084 13976 26140
rect 13912 26080 13976 26084
rect 13992 26140 14056 26144
rect 13992 26084 13996 26140
rect 13996 26084 14052 26140
rect 14052 26084 14056 26140
rect 13992 26080 14056 26084
rect 16752 26140 16816 26144
rect 16752 26084 16756 26140
rect 16756 26084 16812 26140
rect 16812 26084 16816 26140
rect 16752 26080 16816 26084
rect 16832 26140 16896 26144
rect 16832 26084 16836 26140
rect 16836 26084 16892 26140
rect 16892 26084 16896 26140
rect 16832 26080 16896 26084
rect 16912 26140 16976 26144
rect 16912 26084 16916 26140
rect 16916 26084 16972 26140
rect 16972 26084 16976 26140
rect 16912 26080 16976 26084
rect 16992 26140 17056 26144
rect 16992 26084 16996 26140
rect 16996 26084 17052 26140
rect 17052 26084 17056 26140
rect 16992 26080 17056 26084
rect 19752 26140 19816 26144
rect 19752 26084 19756 26140
rect 19756 26084 19812 26140
rect 19812 26084 19816 26140
rect 19752 26080 19816 26084
rect 19832 26140 19896 26144
rect 19832 26084 19836 26140
rect 19836 26084 19892 26140
rect 19892 26084 19896 26140
rect 19832 26080 19896 26084
rect 19912 26140 19976 26144
rect 19912 26084 19916 26140
rect 19916 26084 19972 26140
rect 19972 26084 19976 26140
rect 19912 26080 19976 26084
rect 19992 26140 20056 26144
rect 19992 26084 19996 26140
rect 19996 26084 20052 26140
rect 20052 26084 20056 26140
rect 19992 26080 20056 26084
rect 22752 26140 22816 26144
rect 22752 26084 22756 26140
rect 22756 26084 22812 26140
rect 22812 26084 22816 26140
rect 22752 26080 22816 26084
rect 22832 26140 22896 26144
rect 22832 26084 22836 26140
rect 22836 26084 22892 26140
rect 22892 26084 22896 26140
rect 22832 26080 22896 26084
rect 22912 26140 22976 26144
rect 22912 26084 22916 26140
rect 22916 26084 22972 26140
rect 22972 26084 22976 26140
rect 22912 26080 22976 26084
rect 22992 26140 23056 26144
rect 22992 26084 22996 26140
rect 22996 26084 23052 26140
rect 23052 26084 23056 26140
rect 22992 26080 23056 26084
rect 25752 26140 25816 26144
rect 25752 26084 25756 26140
rect 25756 26084 25812 26140
rect 25812 26084 25816 26140
rect 25752 26080 25816 26084
rect 25832 26140 25896 26144
rect 25832 26084 25836 26140
rect 25836 26084 25892 26140
rect 25892 26084 25896 26140
rect 25832 26080 25896 26084
rect 25912 26140 25976 26144
rect 25912 26084 25916 26140
rect 25916 26084 25972 26140
rect 25972 26084 25976 26140
rect 25912 26080 25976 26084
rect 25992 26140 26056 26144
rect 25992 26084 25996 26140
rect 25996 26084 26052 26140
rect 26052 26084 26056 26140
rect 25992 26080 26056 26084
rect 3252 25596 3316 25600
rect 3252 25540 3256 25596
rect 3256 25540 3312 25596
rect 3312 25540 3316 25596
rect 3252 25536 3316 25540
rect 3332 25596 3396 25600
rect 3332 25540 3336 25596
rect 3336 25540 3392 25596
rect 3392 25540 3396 25596
rect 3332 25536 3396 25540
rect 3412 25596 3476 25600
rect 3412 25540 3416 25596
rect 3416 25540 3472 25596
rect 3472 25540 3476 25596
rect 3412 25536 3476 25540
rect 3492 25596 3556 25600
rect 3492 25540 3496 25596
rect 3496 25540 3552 25596
rect 3552 25540 3556 25596
rect 3492 25536 3556 25540
rect 6252 25596 6316 25600
rect 6252 25540 6256 25596
rect 6256 25540 6312 25596
rect 6312 25540 6316 25596
rect 6252 25536 6316 25540
rect 6332 25596 6396 25600
rect 6332 25540 6336 25596
rect 6336 25540 6392 25596
rect 6392 25540 6396 25596
rect 6332 25536 6396 25540
rect 6412 25596 6476 25600
rect 6412 25540 6416 25596
rect 6416 25540 6472 25596
rect 6472 25540 6476 25596
rect 6412 25536 6476 25540
rect 6492 25596 6556 25600
rect 6492 25540 6496 25596
rect 6496 25540 6552 25596
rect 6552 25540 6556 25596
rect 6492 25536 6556 25540
rect 9252 25596 9316 25600
rect 9252 25540 9256 25596
rect 9256 25540 9312 25596
rect 9312 25540 9316 25596
rect 9252 25536 9316 25540
rect 9332 25596 9396 25600
rect 9332 25540 9336 25596
rect 9336 25540 9392 25596
rect 9392 25540 9396 25596
rect 9332 25536 9396 25540
rect 9412 25596 9476 25600
rect 9412 25540 9416 25596
rect 9416 25540 9472 25596
rect 9472 25540 9476 25596
rect 9412 25536 9476 25540
rect 9492 25596 9556 25600
rect 9492 25540 9496 25596
rect 9496 25540 9552 25596
rect 9552 25540 9556 25596
rect 9492 25536 9556 25540
rect 12252 25596 12316 25600
rect 12252 25540 12256 25596
rect 12256 25540 12312 25596
rect 12312 25540 12316 25596
rect 12252 25536 12316 25540
rect 12332 25596 12396 25600
rect 12332 25540 12336 25596
rect 12336 25540 12392 25596
rect 12392 25540 12396 25596
rect 12332 25536 12396 25540
rect 12412 25596 12476 25600
rect 12412 25540 12416 25596
rect 12416 25540 12472 25596
rect 12472 25540 12476 25596
rect 12412 25536 12476 25540
rect 12492 25596 12556 25600
rect 12492 25540 12496 25596
rect 12496 25540 12552 25596
rect 12552 25540 12556 25596
rect 12492 25536 12556 25540
rect 15252 25596 15316 25600
rect 15252 25540 15256 25596
rect 15256 25540 15312 25596
rect 15312 25540 15316 25596
rect 15252 25536 15316 25540
rect 15332 25596 15396 25600
rect 15332 25540 15336 25596
rect 15336 25540 15392 25596
rect 15392 25540 15396 25596
rect 15332 25536 15396 25540
rect 15412 25596 15476 25600
rect 15412 25540 15416 25596
rect 15416 25540 15472 25596
rect 15472 25540 15476 25596
rect 15412 25536 15476 25540
rect 15492 25596 15556 25600
rect 15492 25540 15496 25596
rect 15496 25540 15552 25596
rect 15552 25540 15556 25596
rect 15492 25536 15556 25540
rect 18252 25596 18316 25600
rect 18252 25540 18256 25596
rect 18256 25540 18312 25596
rect 18312 25540 18316 25596
rect 18252 25536 18316 25540
rect 18332 25596 18396 25600
rect 18332 25540 18336 25596
rect 18336 25540 18392 25596
rect 18392 25540 18396 25596
rect 18332 25536 18396 25540
rect 18412 25596 18476 25600
rect 18412 25540 18416 25596
rect 18416 25540 18472 25596
rect 18472 25540 18476 25596
rect 18412 25536 18476 25540
rect 18492 25596 18556 25600
rect 18492 25540 18496 25596
rect 18496 25540 18552 25596
rect 18552 25540 18556 25596
rect 18492 25536 18556 25540
rect 21252 25596 21316 25600
rect 21252 25540 21256 25596
rect 21256 25540 21312 25596
rect 21312 25540 21316 25596
rect 21252 25536 21316 25540
rect 21332 25596 21396 25600
rect 21332 25540 21336 25596
rect 21336 25540 21392 25596
rect 21392 25540 21396 25596
rect 21332 25536 21396 25540
rect 21412 25596 21476 25600
rect 21412 25540 21416 25596
rect 21416 25540 21472 25596
rect 21472 25540 21476 25596
rect 21412 25536 21476 25540
rect 21492 25596 21556 25600
rect 21492 25540 21496 25596
rect 21496 25540 21552 25596
rect 21552 25540 21556 25596
rect 21492 25536 21556 25540
rect 24252 25596 24316 25600
rect 24252 25540 24256 25596
rect 24256 25540 24312 25596
rect 24312 25540 24316 25596
rect 24252 25536 24316 25540
rect 24332 25596 24396 25600
rect 24332 25540 24336 25596
rect 24336 25540 24392 25596
rect 24392 25540 24396 25596
rect 24332 25536 24396 25540
rect 24412 25596 24476 25600
rect 24412 25540 24416 25596
rect 24416 25540 24472 25596
rect 24472 25540 24476 25596
rect 24412 25536 24476 25540
rect 24492 25596 24556 25600
rect 24492 25540 24496 25596
rect 24496 25540 24552 25596
rect 24552 25540 24556 25596
rect 24492 25536 24556 25540
rect 27252 25596 27316 25600
rect 27252 25540 27256 25596
rect 27256 25540 27312 25596
rect 27312 25540 27316 25596
rect 27252 25536 27316 25540
rect 27332 25596 27396 25600
rect 27332 25540 27336 25596
rect 27336 25540 27392 25596
rect 27392 25540 27396 25596
rect 27332 25536 27396 25540
rect 27412 25596 27476 25600
rect 27412 25540 27416 25596
rect 27416 25540 27472 25596
rect 27472 25540 27476 25596
rect 27412 25536 27476 25540
rect 27492 25596 27556 25600
rect 27492 25540 27496 25596
rect 27496 25540 27552 25596
rect 27552 25540 27556 25596
rect 27492 25536 27556 25540
rect 1752 25052 1816 25056
rect 1752 24996 1756 25052
rect 1756 24996 1812 25052
rect 1812 24996 1816 25052
rect 1752 24992 1816 24996
rect 1832 25052 1896 25056
rect 1832 24996 1836 25052
rect 1836 24996 1892 25052
rect 1892 24996 1896 25052
rect 1832 24992 1896 24996
rect 1912 25052 1976 25056
rect 1912 24996 1916 25052
rect 1916 24996 1972 25052
rect 1972 24996 1976 25052
rect 1912 24992 1976 24996
rect 1992 25052 2056 25056
rect 1992 24996 1996 25052
rect 1996 24996 2052 25052
rect 2052 24996 2056 25052
rect 1992 24992 2056 24996
rect 4752 25052 4816 25056
rect 4752 24996 4756 25052
rect 4756 24996 4812 25052
rect 4812 24996 4816 25052
rect 4752 24992 4816 24996
rect 4832 25052 4896 25056
rect 4832 24996 4836 25052
rect 4836 24996 4892 25052
rect 4892 24996 4896 25052
rect 4832 24992 4896 24996
rect 4912 25052 4976 25056
rect 4912 24996 4916 25052
rect 4916 24996 4972 25052
rect 4972 24996 4976 25052
rect 4912 24992 4976 24996
rect 4992 25052 5056 25056
rect 4992 24996 4996 25052
rect 4996 24996 5052 25052
rect 5052 24996 5056 25052
rect 4992 24992 5056 24996
rect 7752 25052 7816 25056
rect 7752 24996 7756 25052
rect 7756 24996 7812 25052
rect 7812 24996 7816 25052
rect 7752 24992 7816 24996
rect 7832 25052 7896 25056
rect 7832 24996 7836 25052
rect 7836 24996 7892 25052
rect 7892 24996 7896 25052
rect 7832 24992 7896 24996
rect 7912 25052 7976 25056
rect 7912 24996 7916 25052
rect 7916 24996 7972 25052
rect 7972 24996 7976 25052
rect 7912 24992 7976 24996
rect 7992 25052 8056 25056
rect 7992 24996 7996 25052
rect 7996 24996 8052 25052
rect 8052 24996 8056 25052
rect 7992 24992 8056 24996
rect 10752 25052 10816 25056
rect 10752 24996 10756 25052
rect 10756 24996 10812 25052
rect 10812 24996 10816 25052
rect 10752 24992 10816 24996
rect 10832 25052 10896 25056
rect 10832 24996 10836 25052
rect 10836 24996 10892 25052
rect 10892 24996 10896 25052
rect 10832 24992 10896 24996
rect 10912 25052 10976 25056
rect 10912 24996 10916 25052
rect 10916 24996 10972 25052
rect 10972 24996 10976 25052
rect 10912 24992 10976 24996
rect 10992 25052 11056 25056
rect 10992 24996 10996 25052
rect 10996 24996 11052 25052
rect 11052 24996 11056 25052
rect 10992 24992 11056 24996
rect 13752 25052 13816 25056
rect 13752 24996 13756 25052
rect 13756 24996 13812 25052
rect 13812 24996 13816 25052
rect 13752 24992 13816 24996
rect 13832 25052 13896 25056
rect 13832 24996 13836 25052
rect 13836 24996 13892 25052
rect 13892 24996 13896 25052
rect 13832 24992 13896 24996
rect 13912 25052 13976 25056
rect 13912 24996 13916 25052
rect 13916 24996 13972 25052
rect 13972 24996 13976 25052
rect 13912 24992 13976 24996
rect 13992 25052 14056 25056
rect 13992 24996 13996 25052
rect 13996 24996 14052 25052
rect 14052 24996 14056 25052
rect 13992 24992 14056 24996
rect 16752 25052 16816 25056
rect 16752 24996 16756 25052
rect 16756 24996 16812 25052
rect 16812 24996 16816 25052
rect 16752 24992 16816 24996
rect 16832 25052 16896 25056
rect 16832 24996 16836 25052
rect 16836 24996 16892 25052
rect 16892 24996 16896 25052
rect 16832 24992 16896 24996
rect 16912 25052 16976 25056
rect 16912 24996 16916 25052
rect 16916 24996 16972 25052
rect 16972 24996 16976 25052
rect 16912 24992 16976 24996
rect 16992 25052 17056 25056
rect 16992 24996 16996 25052
rect 16996 24996 17052 25052
rect 17052 24996 17056 25052
rect 16992 24992 17056 24996
rect 19752 25052 19816 25056
rect 19752 24996 19756 25052
rect 19756 24996 19812 25052
rect 19812 24996 19816 25052
rect 19752 24992 19816 24996
rect 19832 25052 19896 25056
rect 19832 24996 19836 25052
rect 19836 24996 19892 25052
rect 19892 24996 19896 25052
rect 19832 24992 19896 24996
rect 19912 25052 19976 25056
rect 19912 24996 19916 25052
rect 19916 24996 19972 25052
rect 19972 24996 19976 25052
rect 19912 24992 19976 24996
rect 19992 25052 20056 25056
rect 19992 24996 19996 25052
rect 19996 24996 20052 25052
rect 20052 24996 20056 25052
rect 19992 24992 20056 24996
rect 22752 25052 22816 25056
rect 22752 24996 22756 25052
rect 22756 24996 22812 25052
rect 22812 24996 22816 25052
rect 22752 24992 22816 24996
rect 22832 25052 22896 25056
rect 22832 24996 22836 25052
rect 22836 24996 22892 25052
rect 22892 24996 22896 25052
rect 22832 24992 22896 24996
rect 22912 25052 22976 25056
rect 22912 24996 22916 25052
rect 22916 24996 22972 25052
rect 22972 24996 22976 25052
rect 22912 24992 22976 24996
rect 22992 25052 23056 25056
rect 22992 24996 22996 25052
rect 22996 24996 23052 25052
rect 23052 24996 23056 25052
rect 22992 24992 23056 24996
rect 25752 25052 25816 25056
rect 25752 24996 25756 25052
rect 25756 24996 25812 25052
rect 25812 24996 25816 25052
rect 25752 24992 25816 24996
rect 25832 25052 25896 25056
rect 25832 24996 25836 25052
rect 25836 24996 25892 25052
rect 25892 24996 25896 25052
rect 25832 24992 25896 24996
rect 25912 25052 25976 25056
rect 25912 24996 25916 25052
rect 25916 24996 25972 25052
rect 25972 24996 25976 25052
rect 25912 24992 25976 24996
rect 25992 25052 26056 25056
rect 25992 24996 25996 25052
rect 25996 24996 26052 25052
rect 26052 24996 26056 25052
rect 25992 24992 26056 24996
rect 3252 24508 3316 24512
rect 3252 24452 3256 24508
rect 3256 24452 3312 24508
rect 3312 24452 3316 24508
rect 3252 24448 3316 24452
rect 3332 24508 3396 24512
rect 3332 24452 3336 24508
rect 3336 24452 3392 24508
rect 3392 24452 3396 24508
rect 3332 24448 3396 24452
rect 3412 24508 3476 24512
rect 3412 24452 3416 24508
rect 3416 24452 3472 24508
rect 3472 24452 3476 24508
rect 3412 24448 3476 24452
rect 3492 24508 3556 24512
rect 3492 24452 3496 24508
rect 3496 24452 3552 24508
rect 3552 24452 3556 24508
rect 3492 24448 3556 24452
rect 6252 24508 6316 24512
rect 6252 24452 6256 24508
rect 6256 24452 6312 24508
rect 6312 24452 6316 24508
rect 6252 24448 6316 24452
rect 6332 24508 6396 24512
rect 6332 24452 6336 24508
rect 6336 24452 6392 24508
rect 6392 24452 6396 24508
rect 6332 24448 6396 24452
rect 6412 24508 6476 24512
rect 6412 24452 6416 24508
rect 6416 24452 6472 24508
rect 6472 24452 6476 24508
rect 6412 24448 6476 24452
rect 6492 24508 6556 24512
rect 6492 24452 6496 24508
rect 6496 24452 6552 24508
rect 6552 24452 6556 24508
rect 6492 24448 6556 24452
rect 9252 24508 9316 24512
rect 9252 24452 9256 24508
rect 9256 24452 9312 24508
rect 9312 24452 9316 24508
rect 9252 24448 9316 24452
rect 9332 24508 9396 24512
rect 9332 24452 9336 24508
rect 9336 24452 9392 24508
rect 9392 24452 9396 24508
rect 9332 24448 9396 24452
rect 9412 24508 9476 24512
rect 9412 24452 9416 24508
rect 9416 24452 9472 24508
rect 9472 24452 9476 24508
rect 9412 24448 9476 24452
rect 9492 24508 9556 24512
rect 9492 24452 9496 24508
rect 9496 24452 9552 24508
rect 9552 24452 9556 24508
rect 9492 24448 9556 24452
rect 12252 24508 12316 24512
rect 12252 24452 12256 24508
rect 12256 24452 12312 24508
rect 12312 24452 12316 24508
rect 12252 24448 12316 24452
rect 12332 24508 12396 24512
rect 12332 24452 12336 24508
rect 12336 24452 12392 24508
rect 12392 24452 12396 24508
rect 12332 24448 12396 24452
rect 12412 24508 12476 24512
rect 12412 24452 12416 24508
rect 12416 24452 12472 24508
rect 12472 24452 12476 24508
rect 12412 24448 12476 24452
rect 12492 24508 12556 24512
rect 12492 24452 12496 24508
rect 12496 24452 12552 24508
rect 12552 24452 12556 24508
rect 12492 24448 12556 24452
rect 15252 24508 15316 24512
rect 15252 24452 15256 24508
rect 15256 24452 15312 24508
rect 15312 24452 15316 24508
rect 15252 24448 15316 24452
rect 15332 24508 15396 24512
rect 15332 24452 15336 24508
rect 15336 24452 15392 24508
rect 15392 24452 15396 24508
rect 15332 24448 15396 24452
rect 15412 24508 15476 24512
rect 15412 24452 15416 24508
rect 15416 24452 15472 24508
rect 15472 24452 15476 24508
rect 15412 24448 15476 24452
rect 15492 24508 15556 24512
rect 15492 24452 15496 24508
rect 15496 24452 15552 24508
rect 15552 24452 15556 24508
rect 15492 24448 15556 24452
rect 18252 24508 18316 24512
rect 18252 24452 18256 24508
rect 18256 24452 18312 24508
rect 18312 24452 18316 24508
rect 18252 24448 18316 24452
rect 18332 24508 18396 24512
rect 18332 24452 18336 24508
rect 18336 24452 18392 24508
rect 18392 24452 18396 24508
rect 18332 24448 18396 24452
rect 18412 24508 18476 24512
rect 18412 24452 18416 24508
rect 18416 24452 18472 24508
rect 18472 24452 18476 24508
rect 18412 24448 18476 24452
rect 18492 24508 18556 24512
rect 18492 24452 18496 24508
rect 18496 24452 18552 24508
rect 18552 24452 18556 24508
rect 18492 24448 18556 24452
rect 21252 24508 21316 24512
rect 21252 24452 21256 24508
rect 21256 24452 21312 24508
rect 21312 24452 21316 24508
rect 21252 24448 21316 24452
rect 21332 24508 21396 24512
rect 21332 24452 21336 24508
rect 21336 24452 21392 24508
rect 21392 24452 21396 24508
rect 21332 24448 21396 24452
rect 21412 24508 21476 24512
rect 21412 24452 21416 24508
rect 21416 24452 21472 24508
rect 21472 24452 21476 24508
rect 21412 24448 21476 24452
rect 21492 24508 21556 24512
rect 21492 24452 21496 24508
rect 21496 24452 21552 24508
rect 21552 24452 21556 24508
rect 21492 24448 21556 24452
rect 24252 24508 24316 24512
rect 24252 24452 24256 24508
rect 24256 24452 24312 24508
rect 24312 24452 24316 24508
rect 24252 24448 24316 24452
rect 24332 24508 24396 24512
rect 24332 24452 24336 24508
rect 24336 24452 24392 24508
rect 24392 24452 24396 24508
rect 24332 24448 24396 24452
rect 24412 24508 24476 24512
rect 24412 24452 24416 24508
rect 24416 24452 24472 24508
rect 24472 24452 24476 24508
rect 24412 24448 24476 24452
rect 24492 24508 24556 24512
rect 24492 24452 24496 24508
rect 24496 24452 24552 24508
rect 24552 24452 24556 24508
rect 24492 24448 24556 24452
rect 27252 24508 27316 24512
rect 27252 24452 27256 24508
rect 27256 24452 27312 24508
rect 27312 24452 27316 24508
rect 27252 24448 27316 24452
rect 27332 24508 27396 24512
rect 27332 24452 27336 24508
rect 27336 24452 27392 24508
rect 27392 24452 27396 24508
rect 27332 24448 27396 24452
rect 27412 24508 27476 24512
rect 27412 24452 27416 24508
rect 27416 24452 27472 24508
rect 27472 24452 27476 24508
rect 27412 24448 27476 24452
rect 27492 24508 27556 24512
rect 27492 24452 27496 24508
rect 27496 24452 27552 24508
rect 27552 24452 27556 24508
rect 27492 24448 27556 24452
rect 1752 23964 1816 23968
rect 1752 23908 1756 23964
rect 1756 23908 1812 23964
rect 1812 23908 1816 23964
rect 1752 23904 1816 23908
rect 1832 23964 1896 23968
rect 1832 23908 1836 23964
rect 1836 23908 1892 23964
rect 1892 23908 1896 23964
rect 1832 23904 1896 23908
rect 1912 23964 1976 23968
rect 1912 23908 1916 23964
rect 1916 23908 1972 23964
rect 1972 23908 1976 23964
rect 1912 23904 1976 23908
rect 1992 23964 2056 23968
rect 1992 23908 1996 23964
rect 1996 23908 2052 23964
rect 2052 23908 2056 23964
rect 1992 23904 2056 23908
rect 4752 23964 4816 23968
rect 4752 23908 4756 23964
rect 4756 23908 4812 23964
rect 4812 23908 4816 23964
rect 4752 23904 4816 23908
rect 4832 23964 4896 23968
rect 4832 23908 4836 23964
rect 4836 23908 4892 23964
rect 4892 23908 4896 23964
rect 4832 23904 4896 23908
rect 4912 23964 4976 23968
rect 4912 23908 4916 23964
rect 4916 23908 4972 23964
rect 4972 23908 4976 23964
rect 4912 23904 4976 23908
rect 4992 23964 5056 23968
rect 4992 23908 4996 23964
rect 4996 23908 5052 23964
rect 5052 23908 5056 23964
rect 4992 23904 5056 23908
rect 7752 23964 7816 23968
rect 7752 23908 7756 23964
rect 7756 23908 7812 23964
rect 7812 23908 7816 23964
rect 7752 23904 7816 23908
rect 7832 23964 7896 23968
rect 7832 23908 7836 23964
rect 7836 23908 7892 23964
rect 7892 23908 7896 23964
rect 7832 23904 7896 23908
rect 7912 23964 7976 23968
rect 7912 23908 7916 23964
rect 7916 23908 7972 23964
rect 7972 23908 7976 23964
rect 7912 23904 7976 23908
rect 7992 23964 8056 23968
rect 7992 23908 7996 23964
rect 7996 23908 8052 23964
rect 8052 23908 8056 23964
rect 7992 23904 8056 23908
rect 10752 23964 10816 23968
rect 10752 23908 10756 23964
rect 10756 23908 10812 23964
rect 10812 23908 10816 23964
rect 10752 23904 10816 23908
rect 10832 23964 10896 23968
rect 10832 23908 10836 23964
rect 10836 23908 10892 23964
rect 10892 23908 10896 23964
rect 10832 23904 10896 23908
rect 10912 23964 10976 23968
rect 10912 23908 10916 23964
rect 10916 23908 10972 23964
rect 10972 23908 10976 23964
rect 10912 23904 10976 23908
rect 10992 23964 11056 23968
rect 10992 23908 10996 23964
rect 10996 23908 11052 23964
rect 11052 23908 11056 23964
rect 10992 23904 11056 23908
rect 13752 23964 13816 23968
rect 13752 23908 13756 23964
rect 13756 23908 13812 23964
rect 13812 23908 13816 23964
rect 13752 23904 13816 23908
rect 13832 23964 13896 23968
rect 13832 23908 13836 23964
rect 13836 23908 13892 23964
rect 13892 23908 13896 23964
rect 13832 23904 13896 23908
rect 13912 23964 13976 23968
rect 13912 23908 13916 23964
rect 13916 23908 13972 23964
rect 13972 23908 13976 23964
rect 13912 23904 13976 23908
rect 13992 23964 14056 23968
rect 13992 23908 13996 23964
rect 13996 23908 14052 23964
rect 14052 23908 14056 23964
rect 13992 23904 14056 23908
rect 16752 23964 16816 23968
rect 16752 23908 16756 23964
rect 16756 23908 16812 23964
rect 16812 23908 16816 23964
rect 16752 23904 16816 23908
rect 16832 23964 16896 23968
rect 16832 23908 16836 23964
rect 16836 23908 16892 23964
rect 16892 23908 16896 23964
rect 16832 23904 16896 23908
rect 16912 23964 16976 23968
rect 16912 23908 16916 23964
rect 16916 23908 16972 23964
rect 16972 23908 16976 23964
rect 16912 23904 16976 23908
rect 16992 23964 17056 23968
rect 16992 23908 16996 23964
rect 16996 23908 17052 23964
rect 17052 23908 17056 23964
rect 16992 23904 17056 23908
rect 19752 23964 19816 23968
rect 19752 23908 19756 23964
rect 19756 23908 19812 23964
rect 19812 23908 19816 23964
rect 19752 23904 19816 23908
rect 19832 23964 19896 23968
rect 19832 23908 19836 23964
rect 19836 23908 19892 23964
rect 19892 23908 19896 23964
rect 19832 23904 19896 23908
rect 19912 23964 19976 23968
rect 19912 23908 19916 23964
rect 19916 23908 19972 23964
rect 19972 23908 19976 23964
rect 19912 23904 19976 23908
rect 19992 23964 20056 23968
rect 19992 23908 19996 23964
rect 19996 23908 20052 23964
rect 20052 23908 20056 23964
rect 19992 23904 20056 23908
rect 22752 23964 22816 23968
rect 22752 23908 22756 23964
rect 22756 23908 22812 23964
rect 22812 23908 22816 23964
rect 22752 23904 22816 23908
rect 22832 23964 22896 23968
rect 22832 23908 22836 23964
rect 22836 23908 22892 23964
rect 22892 23908 22896 23964
rect 22832 23904 22896 23908
rect 22912 23964 22976 23968
rect 22912 23908 22916 23964
rect 22916 23908 22972 23964
rect 22972 23908 22976 23964
rect 22912 23904 22976 23908
rect 22992 23964 23056 23968
rect 22992 23908 22996 23964
rect 22996 23908 23052 23964
rect 23052 23908 23056 23964
rect 22992 23904 23056 23908
rect 25752 23964 25816 23968
rect 25752 23908 25756 23964
rect 25756 23908 25812 23964
rect 25812 23908 25816 23964
rect 25752 23904 25816 23908
rect 25832 23964 25896 23968
rect 25832 23908 25836 23964
rect 25836 23908 25892 23964
rect 25892 23908 25896 23964
rect 25832 23904 25896 23908
rect 25912 23964 25976 23968
rect 25912 23908 25916 23964
rect 25916 23908 25972 23964
rect 25972 23908 25976 23964
rect 25912 23904 25976 23908
rect 25992 23964 26056 23968
rect 25992 23908 25996 23964
rect 25996 23908 26052 23964
rect 26052 23908 26056 23964
rect 25992 23904 26056 23908
rect 3252 23420 3316 23424
rect 3252 23364 3256 23420
rect 3256 23364 3312 23420
rect 3312 23364 3316 23420
rect 3252 23360 3316 23364
rect 3332 23420 3396 23424
rect 3332 23364 3336 23420
rect 3336 23364 3392 23420
rect 3392 23364 3396 23420
rect 3332 23360 3396 23364
rect 3412 23420 3476 23424
rect 3412 23364 3416 23420
rect 3416 23364 3472 23420
rect 3472 23364 3476 23420
rect 3412 23360 3476 23364
rect 3492 23420 3556 23424
rect 3492 23364 3496 23420
rect 3496 23364 3552 23420
rect 3552 23364 3556 23420
rect 3492 23360 3556 23364
rect 6252 23420 6316 23424
rect 6252 23364 6256 23420
rect 6256 23364 6312 23420
rect 6312 23364 6316 23420
rect 6252 23360 6316 23364
rect 6332 23420 6396 23424
rect 6332 23364 6336 23420
rect 6336 23364 6392 23420
rect 6392 23364 6396 23420
rect 6332 23360 6396 23364
rect 6412 23420 6476 23424
rect 6412 23364 6416 23420
rect 6416 23364 6472 23420
rect 6472 23364 6476 23420
rect 6412 23360 6476 23364
rect 6492 23420 6556 23424
rect 6492 23364 6496 23420
rect 6496 23364 6552 23420
rect 6552 23364 6556 23420
rect 6492 23360 6556 23364
rect 9252 23420 9316 23424
rect 9252 23364 9256 23420
rect 9256 23364 9312 23420
rect 9312 23364 9316 23420
rect 9252 23360 9316 23364
rect 9332 23420 9396 23424
rect 9332 23364 9336 23420
rect 9336 23364 9392 23420
rect 9392 23364 9396 23420
rect 9332 23360 9396 23364
rect 9412 23420 9476 23424
rect 9412 23364 9416 23420
rect 9416 23364 9472 23420
rect 9472 23364 9476 23420
rect 9412 23360 9476 23364
rect 9492 23420 9556 23424
rect 9492 23364 9496 23420
rect 9496 23364 9552 23420
rect 9552 23364 9556 23420
rect 9492 23360 9556 23364
rect 12252 23420 12316 23424
rect 12252 23364 12256 23420
rect 12256 23364 12312 23420
rect 12312 23364 12316 23420
rect 12252 23360 12316 23364
rect 12332 23420 12396 23424
rect 12332 23364 12336 23420
rect 12336 23364 12392 23420
rect 12392 23364 12396 23420
rect 12332 23360 12396 23364
rect 12412 23420 12476 23424
rect 12412 23364 12416 23420
rect 12416 23364 12472 23420
rect 12472 23364 12476 23420
rect 12412 23360 12476 23364
rect 12492 23420 12556 23424
rect 12492 23364 12496 23420
rect 12496 23364 12552 23420
rect 12552 23364 12556 23420
rect 12492 23360 12556 23364
rect 15252 23420 15316 23424
rect 15252 23364 15256 23420
rect 15256 23364 15312 23420
rect 15312 23364 15316 23420
rect 15252 23360 15316 23364
rect 15332 23420 15396 23424
rect 15332 23364 15336 23420
rect 15336 23364 15392 23420
rect 15392 23364 15396 23420
rect 15332 23360 15396 23364
rect 15412 23420 15476 23424
rect 15412 23364 15416 23420
rect 15416 23364 15472 23420
rect 15472 23364 15476 23420
rect 15412 23360 15476 23364
rect 15492 23420 15556 23424
rect 15492 23364 15496 23420
rect 15496 23364 15552 23420
rect 15552 23364 15556 23420
rect 15492 23360 15556 23364
rect 18252 23420 18316 23424
rect 18252 23364 18256 23420
rect 18256 23364 18312 23420
rect 18312 23364 18316 23420
rect 18252 23360 18316 23364
rect 18332 23420 18396 23424
rect 18332 23364 18336 23420
rect 18336 23364 18392 23420
rect 18392 23364 18396 23420
rect 18332 23360 18396 23364
rect 18412 23420 18476 23424
rect 18412 23364 18416 23420
rect 18416 23364 18472 23420
rect 18472 23364 18476 23420
rect 18412 23360 18476 23364
rect 18492 23420 18556 23424
rect 18492 23364 18496 23420
rect 18496 23364 18552 23420
rect 18552 23364 18556 23420
rect 18492 23360 18556 23364
rect 21252 23420 21316 23424
rect 21252 23364 21256 23420
rect 21256 23364 21312 23420
rect 21312 23364 21316 23420
rect 21252 23360 21316 23364
rect 21332 23420 21396 23424
rect 21332 23364 21336 23420
rect 21336 23364 21392 23420
rect 21392 23364 21396 23420
rect 21332 23360 21396 23364
rect 21412 23420 21476 23424
rect 21412 23364 21416 23420
rect 21416 23364 21472 23420
rect 21472 23364 21476 23420
rect 21412 23360 21476 23364
rect 21492 23420 21556 23424
rect 21492 23364 21496 23420
rect 21496 23364 21552 23420
rect 21552 23364 21556 23420
rect 21492 23360 21556 23364
rect 24252 23420 24316 23424
rect 24252 23364 24256 23420
rect 24256 23364 24312 23420
rect 24312 23364 24316 23420
rect 24252 23360 24316 23364
rect 24332 23420 24396 23424
rect 24332 23364 24336 23420
rect 24336 23364 24392 23420
rect 24392 23364 24396 23420
rect 24332 23360 24396 23364
rect 24412 23420 24476 23424
rect 24412 23364 24416 23420
rect 24416 23364 24472 23420
rect 24472 23364 24476 23420
rect 24412 23360 24476 23364
rect 24492 23420 24556 23424
rect 24492 23364 24496 23420
rect 24496 23364 24552 23420
rect 24552 23364 24556 23420
rect 24492 23360 24556 23364
rect 27252 23420 27316 23424
rect 27252 23364 27256 23420
rect 27256 23364 27312 23420
rect 27312 23364 27316 23420
rect 27252 23360 27316 23364
rect 27332 23420 27396 23424
rect 27332 23364 27336 23420
rect 27336 23364 27392 23420
rect 27392 23364 27396 23420
rect 27332 23360 27396 23364
rect 27412 23420 27476 23424
rect 27412 23364 27416 23420
rect 27416 23364 27472 23420
rect 27472 23364 27476 23420
rect 27412 23360 27476 23364
rect 27492 23420 27556 23424
rect 27492 23364 27496 23420
rect 27496 23364 27552 23420
rect 27552 23364 27556 23420
rect 27492 23360 27556 23364
rect 1752 22876 1816 22880
rect 1752 22820 1756 22876
rect 1756 22820 1812 22876
rect 1812 22820 1816 22876
rect 1752 22816 1816 22820
rect 1832 22876 1896 22880
rect 1832 22820 1836 22876
rect 1836 22820 1892 22876
rect 1892 22820 1896 22876
rect 1832 22816 1896 22820
rect 1912 22876 1976 22880
rect 1912 22820 1916 22876
rect 1916 22820 1972 22876
rect 1972 22820 1976 22876
rect 1912 22816 1976 22820
rect 1992 22876 2056 22880
rect 1992 22820 1996 22876
rect 1996 22820 2052 22876
rect 2052 22820 2056 22876
rect 1992 22816 2056 22820
rect 4752 22876 4816 22880
rect 4752 22820 4756 22876
rect 4756 22820 4812 22876
rect 4812 22820 4816 22876
rect 4752 22816 4816 22820
rect 4832 22876 4896 22880
rect 4832 22820 4836 22876
rect 4836 22820 4892 22876
rect 4892 22820 4896 22876
rect 4832 22816 4896 22820
rect 4912 22876 4976 22880
rect 4912 22820 4916 22876
rect 4916 22820 4972 22876
rect 4972 22820 4976 22876
rect 4912 22816 4976 22820
rect 4992 22876 5056 22880
rect 4992 22820 4996 22876
rect 4996 22820 5052 22876
rect 5052 22820 5056 22876
rect 4992 22816 5056 22820
rect 7752 22876 7816 22880
rect 7752 22820 7756 22876
rect 7756 22820 7812 22876
rect 7812 22820 7816 22876
rect 7752 22816 7816 22820
rect 7832 22876 7896 22880
rect 7832 22820 7836 22876
rect 7836 22820 7892 22876
rect 7892 22820 7896 22876
rect 7832 22816 7896 22820
rect 7912 22876 7976 22880
rect 7912 22820 7916 22876
rect 7916 22820 7972 22876
rect 7972 22820 7976 22876
rect 7912 22816 7976 22820
rect 7992 22876 8056 22880
rect 7992 22820 7996 22876
rect 7996 22820 8052 22876
rect 8052 22820 8056 22876
rect 7992 22816 8056 22820
rect 10752 22876 10816 22880
rect 10752 22820 10756 22876
rect 10756 22820 10812 22876
rect 10812 22820 10816 22876
rect 10752 22816 10816 22820
rect 10832 22876 10896 22880
rect 10832 22820 10836 22876
rect 10836 22820 10892 22876
rect 10892 22820 10896 22876
rect 10832 22816 10896 22820
rect 10912 22876 10976 22880
rect 10912 22820 10916 22876
rect 10916 22820 10972 22876
rect 10972 22820 10976 22876
rect 10912 22816 10976 22820
rect 10992 22876 11056 22880
rect 10992 22820 10996 22876
rect 10996 22820 11052 22876
rect 11052 22820 11056 22876
rect 10992 22816 11056 22820
rect 13752 22876 13816 22880
rect 13752 22820 13756 22876
rect 13756 22820 13812 22876
rect 13812 22820 13816 22876
rect 13752 22816 13816 22820
rect 13832 22876 13896 22880
rect 13832 22820 13836 22876
rect 13836 22820 13892 22876
rect 13892 22820 13896 22876
rect 13832 22816 13896 22820
rect 13912 22876 13976 22880
rect 13912 22820 13916 22876
rect 13916 22820 13972 22876
rect 13972 22820 13976 22876
rect 13912 22816 13976 22820
rect 13992 22876 14056 22880
rect 13992 22820 13996 22876
rect 13996 22820 14052 22876
rect 14052 22820 14056 22876
rect 13992 22816 14056 22820
rect 16752 22876 16816 22880
rect 16752 22820 16756 22876
rect 16756 22820 16812 22876
rect 16812 22820 16816 22876
rect 16752 22816 16816 22820
rect 16832 22876 16896 22880
rect 16832 22820 16836 22876
rect 16836 22820 16892 22876
rect 16892 22820 16896 22876
rect 16832 22816 16896 22820
rect 16912 22876 16976 22880
rect 16912 22820 16916 22876
rect 16916 22820 16972 22876
rect 16972 22820 16976 22876
rect 16912 22816 16976 22820
rect 16992 22876 17056 22880
rect 16992 22820 16996 22876
rect 16996 22820 17052 22876
rect 17052 22820 17056 22876
rect 16992 22816 17056 22820
rect 19752 22876 19816 22880
rect 19752 22820 19756 22876
rect 19756 22820 19812 22876
rect 19812 22820 19816 22876
rect 19752 22816 19816 22820
rect 19832 22876 19896 22880
rect 19832 22820 19836 22876
rect 19836 22820 19892 22876
rect 19892 22820 19896 22876
rect 19832 22816 19896 22820
rect 19912 22876 19976 22880
rect 19912 22820 19916 22876
rect 19916 22820 19972 22876
rect 19972 22820 19976 22876
rect 19912 22816 19976 22820
rect 19992 22876 20056 22880
rect 19992 22820 19996 22876
rect 19996 22820 20052 22876
rect 20052 22820 20056 22876
rect 19992 22816 20056 22820
rect 22752 22876 22816 22880
rect 22752 22820 22756 22876
rect 22756 22820 22812 22876
rect 22812 22820 22816 22876
rect 22752 22816 22816 22820
rect 22832 22876 22896 22880
rect 22832 22820 22836 22876
rect 22836 22820 22892 22876
rect 22892 22820 22896 22876
rect 22832 22816 22896 22820
rect 22912 22876 22976 22880
rect 22912 22820 22916 22876
rect 22916 22820 22972 22876
rect 22972 22820 22976 22876
rect 22912 22816 22976 22820
rect 22992 22876 23056 22880
rect 22992 22820 22996 22876
rect 22996 22820 23052 22876
rect 23052 22820 23056 22876
rect 22992 22816 23056 22820
rect 25752 22876 25816 22880
rect 25752 22820 25756 22876
rect 25756 22820 25812 22876
rect 25812 22820 25816 22876
rect 25752 22816 25816 22820
rect 25832 22876 25896 22880
rect 25832 22820 25836 22876
rect 25836 22820 25892 22876
rect 25892 22820 25896 22876
rect 25832 22816 25896 22820
rect 25912 22876 25976 22880
rect 25912 22820 25916 22876
rect 25916 22820 25972 22876
rect 25972 22820 25976 22876
rect 25912 22816 25976 22820
rect 25992 22876 26056 22880
rect 25992 22820 25996 22876
rect 25996 22820 26052 22876
rect 26052 22820 26056 22876
rect 25992 22816 26056 22820
rect 3252 22332 3316 22336
rect 3252 22276 3256 22332
rect 3256 22276 3312 22332
rect 3312 22276 3316 22332
rect 3252 22272 3316 22276
rect 3332 22332 3396 22336
rect 3332 22276 3336 22332
rect 3336 22276 3392 22332
rect 3392 22276 3396 22332
rect 3332 22272 3396 22276
rect 3412 22332 3476 22336
rect 3412 22276 3416 22332
rect 3416 22276 3472 22332
rect 3472 22276 3476 22332
rect 3412 22272 3476 22276
rect 3492 22332 3556 22336
rect 3492 22276 3496 22332
rect 3496 22276 3552 22332
rect 3552 22276 3556 22332
rect 3492 22272 3556 22276
rect 6252 22332 6316 22336
rect 6252 22276 6256 22332
rect 6256 22276 6312 22332
rect 6312 22276 6316 22332
rect 6252 22272 6316 22276
rect 6332 22332 6396 22336
rect 6332 22276 6336 22332
rect 6336 22276 6392 22332
rect 6392 22276 6396 22332
rect 6332 22272 6396 22276
rect 6412 22332 6476 22336
rect 6412 22276 6416 22332
rect 6416 22276 6472 22332
rect 6472 22276 6476 22332
rect 6412 22272 6476 22276
rect 6492 22332 6556 22336
rect 6492 22276 6496 22332
rect 6496 22276 6552 22332
rect 6552 22276 6556 22332
rect 6492 22272 6556 22276
rect 9252 22332 9316 22336
rect 9252 22276 9256 22332
rect 9256 22276 9312 22332
rect 9312 22276 9316 22332
rect 9252 22272 9316 22276
rect 9332 22332 9396 22336
rect 9332 22276 9336 22332
rect 9336 22276 9392 22332
rect 9392 22276 9396 22332
rect 9332 22272 9396 22276
rect 9412 22332 9476 22336
rect 9412 22276 9416 22332
rect 9416 22276 9472 22332
rect 9472 22276 9476 22332
rect 9412 22272 9476 22276
rect 9492 22332 9556 22336
rect 9492 22276 9496 22332
rect 9496 22276 9552 22332
rect 9552 22276 9556 22332
rect 9492 22272 9556 22276
rect 12252 22332 12316 22336
rect 12252 22276 12256 22332
rect 12256 22276 12312 22332
rect 12312 22276 12316 22332
rect 12252 22272 12316 22276
rect 12332 22332 12396 22336
rect 12332 22276 12336 22332
rect 12336 22276 12392 22332
rect 12392 22276 12396 22332
rect 12332 22272 12396 22276
rect 12412 22332 12476 22336
rect 12412 22276 12416 22332
rect 12416 22276 12472 22332
rect 12472 22276 12476 22332
rect 12412 22272 12476 22276
rect 12492 22332 12556 22336
rect 12492 22276 12496 22332
rect 12496 22276 12552 22332
rect 12552 22276 12556 22332
rect 12492 22272 12556 22276
rect 15252 22332 15316 22336
rect 15252 22276 15256 22332
rect 15256 22276 15312 22332
rect 15312 22276 15316 22332
rect 15252 22272 15316 22276
rect 15332 22332 15396 22336
rect 15332 22276 15336 22332
rect 15336 22276 15392 22332
rect 15392 22276 15396 22332
rect 15332 22272 15396 22276
rect 15412 22332 15476 22336
rect 15412 22276 15416 22332
rect 15416 22276 15472 22332
rect 15472 22276 15476 22332
rect 15412 22272 15476 22276
rect 15492 22332 15556 22336
rect 15492 22276 15496 22332
rect 15496 22276 15552 22332
rect 15552 22276 15556 22332
rect 15492 22272 15556 22276
rect 18252 22332 18316 22336
rect 18252 22276 18256 22332
rect 18256 22276 18312 22332
rect 18312 22276 18316 22332
rect 18252 22272 18316 22276
rect 18332 22332 18396 22336
rect 18332 22276 18336 22332
rect 18336 22276 18392 22332
rect 18392 22276 18396 22332
rect 18332 22272 18396 22276
rect 18412 22332 18476 22336
rect 18412 22276 18416 22332
rect 18416 22276 18472 22332
rect 18472 22276 18476 22332
rect 18412 22272 18476 22276
rect 18492 22332 18556 22336
rect 18492 22276 18496 22332
rect 18496 22276 18552 22332
rect 18552 22276 18556 22332
rect 18492 22272 18556 22276
rect 21252 22332 21316 22336
rect 21252 22276 21256 22332
rect 21256 22276 21312 22332
rect 21312 22276 21316 22332
rect 21252 22272 21316 22276
rect 21332 22332 21396 22336
rect 21332 22276 21336 22332
rect 21336 22276 21392 22332
rect 21392 22276 21396 22332
rect 21332 22272 21396 22276
rect 21412 22332 21476 22336
rect 21412 22276 21416 22332
rect 21416 22276 21472 22332
rect 21472 22276 21476 22332
rect 21412 22272 21476 22276
rect 21492 22332 21556 22336
rect 21492 22276 21496 22332
rect 21496 22276 21552 22332
rect 21552 22276 21556 22332
rect 21492 22272 21556 22276
rect 24252 22332 24316 22336
rect 24252 22276 24256 22332
rect 24256 22276 24312 22332
rect 24312 22276 24316 22332
rect 24252 22272 24316 22276
rect 24332 22332 24396 22336
rect 24332 22276 24336 22332
rect 24336 22276 24392 22332
rect 24392 22276 24396 22332
rect 24332 22272 24396 22276
rect 24412 22332 24476 22336
rect 24412 22276 24416 22332
rect 24416 22276 24472 22332
rect 24472 22276 24476 22332
rect 24412 22272 24476 22276
rect 24492 22332 24556 22336
rect 24492 22276 24496 22332
rect 24496 22276 24552 22332
rect 24552 22276 24556 22332
rect 24492 22272 24556 22276
rect 27252 22332 27316 22336
rect 27252 22276 27256 22332
rect 27256 22276 27312 22332
rect 27312 22276 27316 22332
rect 27252 22272 27316 22276
rect 27332 22332 27396 22336
rect 27332 22276 27336 22332
rect 27336 22276 27392 22332
rect 27392 22276 27396 22332
rect 27332 22272 27396 22276
rect 27412 22332 27476 22336
rect 27412 22276 27416 22332
rect 27416 22276 27472 22332
rect 27472 22276 27476 22332
rect 27412 22272 27476 22276
rect 27492 22332 27556 22336
rect 27492 22276 27496 22332
rect 27496 22276 27552 22332
rect 27552 22276 27556 22332
rect 27492 22272 27556 22276
rect 1752 21788 1816 21792
rect 1752 21732 1756 21788
rect 1756 21732 1812 21788
rect 1812 21732 1816 21788
rect 1752 21728 1816 21732
rect 1832 21788 1896 21792
rect 1832 21732 1836 21788
rect 1836 21732 1892 21788
rect 1892 21732 1896 21788
rect 1832 21728 1896 21732
rect 1912 21788 1976 21792
rect 1912 21732 1916 21788
rect 1916 21732 1972 21788
rect 1972 21732 1976 21788
rect 1912 21728 1976 21732
rect 1992 21788 2056 21792
rect 1992 21732 1996 21788
rect 1996 21732 2052 21788
rect 2052 21732 2056 21788
rect 1992 21728 2056 21732
rect 4752 21788 4816 21792
rect 4752 21732 4756 21788
rect 4756 21732 4812 21788
rect 4812 21732 4816 21788
rect 4752 21728 4816 21732
rect 4832 21788 4896 21792
rect 4832 21732 4836 21788
rect 4836 21732 4892 21788
rect 4892 21732 4896 21788
rect 4832 21728 4896 21732
rect 4912 21788 4976 21792
rect 4912 21732 4916 21788
rect 4916 21732 4972 21788
rect 4972 21732 4976 21788
rect 4912 21728 4976 21732
rect 4992 21788 5056 21792
rect 4992 21732 4996 21788
rect 4996 21732 5052 21788
rect 5052 21732 5056 21788
rect 4992 21728 5056 21732
rect 7752 21788 7816 21792
rect 7752 21732 7756 21788
rect 7756 21732 7812 21788
rect 7812 21732 7816 21788
rect 7752 21728 7816 21732
rect 7832 21788 7896 21792
rect 7832 21732 7836 21788
rect 7836 21732 7892 21788
rect 7892 21732 7896 21788
rect 7832 21728 7896 21732
rect 7912 21788 7976 21792
rect 7912 21732 7916 21788
rect 7916 21732 7972 21788
rect 7972 21732 7976 21788
rect 7912 21728 7976 21732
rect 7992 21788 8056 21792
rect 7992 21732 7996 21788
rect 7996 21732 8052 21788
rect 8052 21732 8056 21788
rect 7992 21728 8056 21732
rect 10752 21788 10816 21792
rect 10752 21732 10756 21788
rect 10756 21732 10812 21788
rect 10812 21732 10816 21788
rect 10752 21728 10816 21732
rect 10832 21788 10896 21792
rect 10832 21732 10836 21788
rect 10836 21732 10892 21788
rect 10892 21732 10896 21788
rect 10832 21728 10896 21732
rect 10912 21788 10976 21792
rect 10912 21732 10916 21788
rect 10916 21732 10972 21788
rect 10972 21732 10976 21788
rect 10912 21728 10976 21732
rect 10992 21788 11056 21792
rect 10992 21732 10996 21788
rect 10996 21732 11052 21788
rect 11052 21732 11056 21788
rect 10992 21728 11056 21732
rect 13752 21788 13816 21792
rect 13752 21732 13756 21788
rect 13756 21732 13812 21788
rect 13812 21732 13816 21788
rect 13752 21728 13816 21732
rect 13832 21788 13896 21792
rect 13832 21732 13836 21788
rect 13836 21732 13892 21788
rect 13892 21732 13896 21788
rect 13832 21728 13896 21732
rect 13912 21788 13976 21792
rect 13912 21732 13916 21788
rect 13916 21732 13972 21788
rect 13972 21732 13976 21788
rect 13912 21728 13976 21732
rect 13992 21788 14056 21792
rect 13992 21732 13996 21788
rect 13996 21732 14052 21788
rect 14052 21732 14056 21788
rect 13992 21728 14056 21732
rect 16752 21788 16816 21792
rect 16752 21732 16756 21788
rect 16756 21732 16812 21788
rect 16812 21732 16816 21788
rect 16752 21728 16816 21732
rect 16832 21788 16896 21792
rect 16832 21732 16836 21788
rect 16836 21732 16892 21788
rect 16892 21732 16896 21788
rect 16832 21728 16896 21732
rect 16912 21788 16976 21792
rect 16912 21732 16916 21788
rect 16916 21732 16972 21788
rect 16972 21732 16976 21788
rect 16912 21728 16976 21732
rect 16992 21788 17056 21792
rect 16992 21732 16996 21788
rect 16996 21732 17052 21788
rect 17052 21732 17056 21788
rect 16992 21728 17056 21732
rect 19752 21788 19816 21792
rect 19752 21732 19756 21788
rect 19756 21732 19812 21788
rect 19812 21732 19816 21788
rect 19752 21728 19816 21732
rect 19832 21788 19896 21792
rect 19832 21732 19836 21788
rect 19836 21732 19892 21788
rect 19892 21732 19896 21788
rect 19832 21728 19896 21732
rect 19912 21788 19976 21792
rect 19912 21732 19916 21788
rect 19916 21732 19972 21788
rect 19972 21732 19976 21788
rect 19912 21728 19976 21732
rect 19992 21788 20056 21792
rect 19992 21732 19996 21788
rect 19996 21732 20052 21788
rect 20052 21732 20056 21788
rect 19992 21728 20056 21732
rect 22752 21788 22816 21792
rect 22752 21732 22756 21788
rect 22756 21732 22812 21788
rect 22812 21732 22816 21788
rect 22752 21728 22816 21732
rect 22832 21788 22896 21792
rect 22832 21732 22836 21788
rect 22836 21732 22892 21788
rect 22892 21732 22896 21788
rect 22832 21728 22896 21732
rect 22912 21788 22976 21792
rect 22912 21732 22916 21788
rect 22916 21732 22972 21788
rect 22972 21732 22976 21788
rect 22912 21728 22976 21732
rect 22992 21788 23056 21792
rect 22992 21732 22996 21788
rect 22996 21732 23052 21788
rect 23052 21732 23056 21788
rect 22992 21728 23056 21732
rect 25752 21788 25816 21792
rect 25752 21732 25756 21788
rect 25756 21732 25812 21788
rect 25812 21732 25816 21788
rect 25752 21728 25816 21732
rect 25832 21788 25896 21792
rect 25832 21732 25836 21788
rect 25836 21732 25892 21788
rect 25892 21732 25896 21788
rect 25832 21728 25896 21732
rect 25912 21788 25976 21792
rect 25912 21732 25916 21788
rect 25916 21732 25972 21788
rect 25972 21732 25976 21788
rect 25912 21728 25976 21732
rect 25992 21788 26056 21792
rect 25992 21732 25996 21788
rect 25996 21732 26052 21788
rect 26052 21732 26056 21788
rect 25992 21728 26056 21732
rect 3252 21244 3316 21248
rect 3252 21188 3256 21244
rect 3256 21188 3312 21244
rect 3312 21188 3316 21244
rect 3252 21184 3316 21188
rect 3332 21244 3396 21248
rect 3332 21188 3336 21244
rect 3336 21188 3392 21244
rect 3392 21188 3396 21244
rect 3332 21184 3396 21188
rect 3412 21244 3476 21248
rect 3412 21188 3416 21244
rect 3416 21188 3472 21244
rect 3472 21188 3476 21244
rect 3412 21184 3476 21188
rect 3492 21244 3556 21248
rect 3492 21188 3496 21244
rect 3496 21188 3552 21244
rect 3552 21188 3556 21244
rect 3492 21184 3556 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 6412 21244 6476 21248
rect 6412 21188 6416 21244
rect 6416 21188 6472 21244
rect 6472 21188 6476 21244
rect 6412 21184 6476 21188
rect 6492 21244 6556 21248
rect 6492 21188 6496 21244
rect 6496 21188 6552 21244
rect 6552 21188 6556 21244
rect 6492 21184 6556 21188
rect 9252 21244 9316 21248
rect 9252 21188 9256 21244
rect 9256 21188 9312 21244
rect 9312 21188 9316 21244
rect 9252 21184 9316 21188
rect 9332 21244 9396 21248
rect 9332 21188 9336 21244
rect 9336 21188 9392 21244
rect 9392 21188 9396 21244
rect 9332 21184 9396 21188
rect 9412 21244 9476 21248
rect 9412 21188 9416 21244
rect 9416 21188 9472 21244
rect 9472 21188 9476 21244
rect 9412 21184 9476 21188
rect 9492 21244 9556 21248
rect 9492 21188 9496 21244
rect 9496 21188 9552 21244
rect 9552 21188 9556 21244
rect 9492 21184 9556 21188
rect 12252 21244 12316 21248
rect 12252 21188 12256 21244
rect 12256 21188 12312 21244
rect 12312 21188 12316 21244
rect 12252 21184 12316 21188
rect 12332 21244 12396 21248
rect 12332 21188 12336 21244
rect 12336 21188 12392 21244
rect 12392 21188 12396 21244
rect 12332 21184 12396 21188
rect 12412 21244 12476 21248
rect 12412 21188 12416 21244
rect 12416 21188 12472 21244
rect 12472 21188 12476 21244
rect 12412 21184 12476 21188
rect 12492 21244 12556 21248
rect 12492 21188 12496 21244
rect 12496 21188 12552 21244
rect 12552 21188 12556 21244
rect 12492 21184 12556 21188
rect 15252 21244 15316 21248
rect 15252 21188 15256 21244
rect 15256 21188 15312 21244
rect 15312 21188 15316 21244
rect 15252 21184 15316 21188
rect 15332 21244 15396 21248
rect 15332 21188 15336 21244
rect 15336 21188 15392 21244
rect 15392 21188 15396 21244
rect 15332 21184 15396 21188
rect 15412 21244 15476 21248
rect 15412 21188 15416 21244
rect 15416 21188 15472 21244
rect 15472 21188 15476 21244
rect 15412 21184 15476 21188
rect 15492 21244 15556 21248
rect 15492 21188 15496 21244
rect 15496 21188 15552 21244
rect 15552 21188 15556 21244
rect 15492 21184 15556 21188
rect 18252 21244 18316 21248
rect 18252 21188 18256 21244
rect 18256 21188 18312 21244
rect 18312 21188 18316 21244
rect 18252 21184 18316 21188
rect 18332 21244 18396 21248
rect 18332 21188 18336 21244
rect 18336 21188 18392 21244
rect 18392 21188 18396 21244
rect 18332 21184 18396 21188
rect 18412 21244 18476 21248
rect 18412 21188 18416 21244
rect 18416 21188 18472 21244
rect 18472 21188 18476 21244
rect 18412 21184 18476 21188
rect 18492 21244 18556 21248
rect 18492 21188 18496 21244
rect 18496 21188 18552 21244
rect 18552 21188 18556 21244
rect 18492 21184 18556 21188
rect 21252 21244 21316 21248
rect 21252 21188 21256 21244
rect 21256 21188 21312 21244
rect 21312 21188 21316 21244
rect 21252 21184 21316 21188
rect 21332 21244 21396 21248
rect 21332 21188 21336 21244
rect 21336 21188 21392 21244
rect 21392 21188 21396 21244
rect 21332 21184 21396 21188
rect 21412 21244 21476 21248
rect 21412 21188 21416 21244
rect 21416 21188 21472 21244
rect 21472 21188 21476 21244
rect 21412 21184 21476 21188
rect 21492 21244 21556 21248
rect 21492 21188 21496 21244
rect 21496 21188 21552 21244
rect 21552 21188 21556 21244
rect 21492 21184 21556 21188
rect 24252 21244 24316 21248
rect 24252 21188 24256 21244
rect 24256 21188 24312 21244
rect 24312 21188 24316 21244
rect 24252 21184 24316 21188
rect 24332 21244 24396 21248
rect 24332 21188 24336 21244
rect 24336 21188 24392 21244
rect 24392 21188 24396 21244
rect 24332 21184 24396 21188
rect 24412 21244 24476 21248
rect 24412 21188 24416 21244
rect 24416 21188 24472 21244
rect 24472 21188 24476 21244
rect 24412 21184 24476 21188
rect 24492 21244 24556 21248
rect 24492 21188 24496 21244
rect 24496 21188 24552 21244
rect 24552 21188 24556 21244
rect 24492 21184 24556 21188
rect 27252 21244 27316 21248
rect 27252 21188 27256 21244
rect 27256 21188 27312 21244
rect 27312 21188 27316 21244
rect 27252 21184 27316 21188
rect 27332 21244 27396 21248
rect 27332 21188 27336 21244
rect 27336 21188 27392 21244
rect 27392 21188 27396 21244
rect 27332 21184 27396 21188
rect 27412 21244 27476 21248
rect 27412 21188 27416 21244
rect 27416 21188 27472 21244
rect 27472 21188 27476 21244
rect 27412 21184 27476 21188
rect 27492 21244 27556 21248
rect 27492 21188 27496 21244
rect 27496 21188 27552 21244
rect 27552 21188 27556 21244
rect 27492 21184 27556 21188
rect 1752 20700 1816 20704
rect 1752 20644 1756 20700
rect 1756 20644 1812 20700
rect 1812 20644 1816 20700
rect 1752 20640 1816 20644
rect 1832 20700 1896 20704
rect 1832 20644 1836 20700
rect 1836 20644 1892 20700
rect 1892 20644 1896 20700
rect 1832 20640 1896 20644
rect 1912 20700 1976 20704
rect 1912 20644 1916 20700
rect 1916 20644 1972 20700
rect 1972 20644 1976 20700
rect 1912 20640 1976 20644
rect 1992 20700 2056 20704
rect 1992 20644 1996 20700
rect 1996 20644 2052 20700
rect 2052 20644 2056 20700
rect 1992 20640 2056 20644
rect 4752 20700 4816 20704
rect 4752 20644 4756 20700
rect 4756 20644 4812 20700
rect 4812 20644 4816 20700
rect 4752 20640 4816 20644
rect 4832 20700 4896 20704
rect 4832 20644 4836 20700
rect 4836 20644 4892 20700
rect 4892 20644 4896 20700
rect 4832 20640 4896 20644
rect 4912 20700 4976 20704
rect 4912 20644 4916 20700
rect 4916 20644 4972 20700
rect 4972 20644 4976 20700
rect 4912 20640 4976 20644
rect 4992 20700 5056 20704
rect 4992 20644 4996 20700
rect 4996 20644 5052 20700
rect 5052 20644 5056 20700
rect 4992 20640 5056 20644
rect 7752 20700 7816 20704
rect 7752 20644 7756 20700
rect 7756 20644 7812 20700
rect 7812 20644 7816 20700
rect 7752 20640 7816 20644
rect 7832 20700 7896 20704
rect 7832 20644 7836 20700
rect 7836 20644 7892 20700
rect 7892 20644 7896 20700
rect 7832 20640 7896 20644
rect 7912 20700 7976 20704
rect 7912 20644 7916 20700
rect 7916 20644 7972 20700
rect 7972 20644 7976 20700
rect 7912 20640 7976 20644
rect 7992 20700 8056 20704
rect 7992 20644 7996 20700
rect 7996 20644 8052 20700
rect 8052 20644 8056 20700
rect 7992 20640 8056 20644
rect 10752 20700 10816 20704
rect 10752 20644 10756 20700
rect 10756 20644 10812 20700
rect 10812 20644 10816 20700
rect 10752 20640 10816 20644
rect 10832 20700 10896 20704
rect 10832 20644 10836 20700
rect 10836 20644 10892 20700
rect 10892 20644 10896 20700
rect 10832 20640 10896 20644
rect 10912 20700 10976 20704
rect 10912 20644 10916 20700
rect 10916 20644 10972 20700
rect 10972 20644 10976 20700
rect 10912 20640 10976 20644
rect 10992 20700 11056 20704
rect 10992 20644 10996 20700
rect 10996 20644 11052 20700
rect 11052 20644 11056 20700
rect 10992 20640 11056 20644
rect 13752 20700 13816 20704
rect 13752 20644 13756 20700
rect 13756 20644 13812 20700
rect 13812 20644 13816 20700
rect 13752 20640 13816 20644
rect 13832 20700 13896 20704
rect 13832 20644 13836 20700
rect 13836 20644 13892 20700
rect 13892 20644 13896 20700
rect 13832 20640 13896 20644
rect 13912 20700 13976 20704
rect 13912 20644 13916 20700
rect 13916 20644 13972 20700
rect 13972 20644 13976 20700
rect 13912 20640 13976 20644
rect 13992 20700 14056 20704
rect 13992 20644 13996 20700
rect 13996 20644 14052 20700
rect 14052 20644 14056 20700
rect 13992 20640 14056 20644
rect 16752 20700 16816 20704
rect 16752 20644 16756 20700
rect 16756 20644 16812 20700
rect 16812 20644 16816 20700
rect 16752 20640 16816 20644
rect 16832 20700 16896 20704
rect 16832 20644 16836 20700
rect 16836 20644 16892 20700
rect 16892 20644 16896 20700
rect 16832 20640 16896 20644
rect 16912 20700 16976 20704
rect 16912 20644 16916 20700
rect 16916 20644 16972 20700
rect 16972 20644 16976 20700
rect 16912 20640 16976 20644
rect 16992 20700 17056 20704
rect 16992 20644 16996 20700
rect 16996 20644 17052 20700
rect 17052 20644 17056 20700
rect 16992 20640 17056 20644
rect 19752 20700 19816 20704
rect 19752 20644 19756 20700
rect 19756 20644 19812 20700
rect 19812 20644 19816 20700
rect 19752 20640 19816 20644
rect 19832 20700 19896 20704
rect 19832 20644 19836 20700
rect 19836 20644 19892 20700
rect 19892 20644 19896 20700
rect 19832 20640 19896 20644
rect 19912 20700 19976 20704
rect 19912 20644 19916 20700
rect 19916 20644 19972 20700
rect 19972 20644 19976 20700
rect 19912 20640 19976 20644
rect 19992 20700 20056 20704
rect 19992 20644 19996 20700
rect 19996 20644 20052 20700
rect 20052 20644 20056 20700
rect 19992 20640 20056 20644
rect 22752 20700 22816 20704
rect 22752 20644 22756 20700
rect 22756 20644 22812 20700
rect 22812 20644 22816 20700
rect 22752 20640 22816 20644
rect 22832 20700 22896 20704
rect 22832 20644 22836 20700
rect 22836 20644 22892 20700
rect 22892 20644 22896 20700
rect 22832 20640 22896 20644
rect 22912 20700 22976 20704
rect 22912 20644 22916 20700
rect 22916 20644 22972 20700
rect 22972 20644 22976 20700
rect 22912 20640 22976 20644
rect 22992 20700 23056 20704
rect 22992 20644 22996 20700
rect 22996 20644 23052 20700
rect 23052 20644 23056 20700
rect 22992 20640 23056 20644
rect 25752 20700 25816 20704
rect 25752 20644 25756 20700
rect 25756 20644 25812 20700
rect 25812 20644 25816 20700
rect 25752 20640 25816 20644
rect 25832 20700 25896 20704
rect 25832 20644 25836 20700
rect 25836 20644 25892 20700
rect 25892 20644 25896 20700
rect 25832 20640 25896 20644
rect 25912 20700 25976 20704
rect 25912 20644 25916 20700
rect 25916 20644 25972 20700
rect 25972 20644 25976 20700
rect 25912 20640 25976 20644
rect 25992 20700 26056 20704
rect 25992 20644 25996 20700
rect 25996 20644 26052 20700
rect 26052 20644 26056 20700
rect 25992 20640 26056 20644
rect 3252 20156 3316 20160
rect 3252 20100 3256 20156
rect 3256 20100 3312 20156
rect 3312 20100 3316 20156
rect 3252 20096 3316 20100
rect 3332 20156 3396 20160
rect 3332 20100 3336 20156
rect 3336 20100 3392 20156
rect 3392 20100 3396 20156
rect 3332 20096 3396 20100
rect 3412 20156 3476 20160
rect 3412 20100 3416 20156
rect 3416 20100 3472 20156
rect 3472 20100 3476 20156
rect 3412 20096 3476 20100
rect 3492 20156 3556 20160
rect 3492 20100 3496 20156
rect 3496 20100 3552 20156
rect 3552 20100 3556 20156
rect 3492 20096 3556 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 6412 20156 6476 20160
rect 6412 20100 6416 20156
rect 6416 20100 6472 20156
rect 6472 20100 6476 20156
rect 6412 20096 6476 20100
rect 6492 20156 6556 20160
rect 6492 20100 6496 20156
rect 6496 20100 6552 20156
rect 6552 20100 6556 20156
rect 6492 20096 6556 20100
rect 9252 20156 9316 20160
rect 9252 20100 9256 20156
rect 9256 20100 9312 20156
rect 9312 20100 9316 20156
rect 9252 20096 9316 20100
rect 9332 20156 9396 20160
rect 9332 20100 9336 20156
rect 9336 20100 9392 20156
rect 9392 20100 9396 20156
rect 9332 20096 9396 20100
rect 9412 20156 9476 20160
rect 9412 20100 9416 20156
rect 9416 20100 9472 20156
rect 9472 20100 9476 20156
rect 9412 20096 9476 20100
rect 9492 20156 9556 20160
rect 9492 20100 9496 20156
rect 9496 20100 9552 20156
rect 9552 20100 9556 20156
rect 9492 20096 9556 20100
rect 12252 20156 12316 20160
rect 12252 20100 12256 20156
rect 12256 20100 12312 20156
rect 12312 20100 12316 20156
rect 12252 20096 12316 20100
rect 12332 20156 12396 20160
rect 12332 20100 12336 20156
rect 12336 20100 12392 20156
rect 12392 20100 12396 20156
rect 12332 20096 12396 20100
rect 12412 20156 12476 20160
rect 12412 20100 12416 20156
rect 12416 20100 12472 20156
rect 12472 20100 12476 20156
rect 12412 20096 12476 20100
rect 12492 20156 12556 20160
rect 12492 20100 12496 20156
rect 12496 20100 12552 20156
rect 12552 20100 12556 20156
rect 12492 20096 12556 20100
rect 15252 20156 15316 20160
rect 15252 20100 15256 20156
rect 15256 20100 15312 20156
rect 15312 20100 15316 20156
rect 15252 20096 15316 20100
rect 15332 20156 15396 20160
rect 15332 20100 15336 20156
rect 15336 20100 15392 20156
rect 15392 20100 15396 20156
rect 15332 20096 15396 20100
rect 15412 20156 15476 20160
rect 15412 20100 15416 20156
rect 15416 20100 15472 20156
rect 15472 20100 15476 20156
rect 15412 20096 15476 20100
rect 15492 20156 15556 20160
rect 15492 20100 15496 20156
rect 15496 20100 15552 20156
rect 15552 20100 15556 20156
rect 15492 20096 15556 20100
rect 18252 20156 18316 20160
rect 18252 20100 18256 20156
rect 18256 20100 18312 20156
rect 18312 20100 18316 20156
rect 18252 20096 18316 20100
rect 18332 20156 18396 20160
rect 18332 20100 18336 20156
rect 18336 20100 18392 20156
rect 18392 20100 18396 20156
rect 18332 20096 18396 20100
rect 18412 20156 18476 20160
rect 18412 20100 18416 20156
rect 18416 20100 18472 20156
rect 18472 20100 18476 20156
rect 18412 20096 18476 20100
rect 18492 20156 18556 20160
rect 18492 20100 18496 20156
rect 18496 20100 18552 20156
rect 18552 20100 18556 20156
rect 18492 20096 18556 20100
rect 21252 20156 21316 20160
rect 21252 20100 21256 20156
rect 21256 20100 21312 20156
rect 21312 20100 21316 20156
rect 21252 20096 21316 20100
rect 21332 20156 21396 20160
rect 21332 20100 21336 20156
rect 21336 20100 21392 20156
rect 21392 20100 21396 20156
rect 21332 20096 21396 20100
rect 21412 20156 21476 20160
rect 21412 20100 21416 20156
rect 21416 20100 21472 20156
rect 21472 20100 21476 20156
rect 21412 20096 21476 20100
rect 21492 20156 21556 20160
rect 21492 20100 21496 20156
rect 21496 20100 21552 20156
rect 21552 20100 21556 20156
rect 21492 20096 21556 20100
rect 24252 20156 24316 20160
rect 24252 20100 24256 20156
rect 24256 20100 24312 20156
rect 24312 20100 24316 20156
rect 24252 20096 24316 20100
rect 24332 20156 24396 20160
rect 24332 20100 24336 20156
rect 24336 20100 24392 20156
rect 24392 20100 24396 20156
rect 24332 20096 24396 20100
rect 24412 20156 24476 20160
rect 24412 20100 24416 20156
rect 24416 20100 24472 20156
rect 24472 20100 24476 20156
rect 24412 20096 24476 20100
rect 24492 20156 24556 20160
rect 24492 20100 24496 20156
rect 24496 20100 24552 20156
rect 24552 20100 24556 20156
rect 24492 20096 24556 20100
rect 27252 20156 27316 20160
rect 27252 20100 27256 20156
rect 27256 20100 27312 20156
rect 27312 20100 27316 20156
rect 27252 20096 27316 20100
rect 27332 20156 27396 20160
rect 27332 20100 27336 20156
rect 27336 20100 27392 20156
rect 27392 20100 27396 20156
rect 27332 20096 27396 20100
rect 27412 20156 27476 20160
rect 27412 20100 27416 20156
rect 27416 20100 27472 20156
rect 27472 20100 27476 20156
rect 27412 20096 27476 20100
rect 27492 20156 27556 20160
rect 27492 20100 27496 20156
rect 27496 20100 27552 20156
rect 27552 20100 27556 20156
rect 27492 20096 27556 20100
rect 1752 19612 1816 19616
rect 1752 19556 1756 19612
rect 1756 19556 1812 19612
rect 1812 19556 1816 19612
rect 1752 19552 1816 19556
rect 1832 19612 1896 19616
rect 1832 19556 1836 19612
rect 1836 19556 1892 19612
rect 1892 19556 1896 19612
rect 1832 19552 1896 19556
rect 1912 19612 1976 19616
rect 1912 19556 1916 19612
rect 1916 19556 1972 19612
rect 1972 19556 1976 19612
rect 1912 19552 1976 19556
rect 1992 19612 2056 19616
rect 1992 19556 1996 19612
rect 1996 19556 2052 19612
rect 2052 19556 2056 19612
rect 1992 19552 2056 19556
rect 4752 19612 4816 19616
rect 4752 19556 4756 19612
rect 4756 19556 4812 19612
rect 4812 19556 4816 19612
rect 4752 19552 4816 19556
rect 4832 19612 4896 19616
rect 4832 19556 4836 19612
rect 4836 19556 4892 19612
rect 4892 19556 4896 19612
rect 4832 19552 4896 19556
rect 4912 19612 4976 19616
rect 4912 19556 4916 19612
rect 4916 19556 4972 19612
rect 4972 19556 4976 19612
rect 4912 19552 4976 19556
rect 4992 19612 5056 19616
rect 4992 19556 4996 19612
rect 4996 19556 5052 19612
rect 5052 19556 5056 19612
rect 4992 19552 5056 19556
rect 7752 19612 7816 19616
rect 7752 19556 7756 19612
rect 7756 19556 7812 19612
rect 7812 19556 7816 19612
rect 7752 19552 7816 19556
rect 7832 19612 7896 19616
rect 7832 19556 7836 19612
rect 7836 19556 7892 19612
rect 7892 19556 7896 19612
rect 7832 19552 7896 19556
rect 7912 19612 7976 19616
rect 7912 19556 7916 19612
rect 7916 19556 7972 19612
rect 7972 19556 7976 19612
rect 7912 19552 7976 19556
rect 7992 19612 8056 19616
rect 7992 19556 7996 19612
rect 7996 19556 8052 19612
rect 8052 19556 8056 19612
rect 7992 19552 8056 19556
rect 10752 19612 10816 19616
rect 10752 19556 10756 19612
rect 10756 19556 10812 19612
rect 10812 19556 10816 19612
rect 10752 19552 10816 19556
rect 10832 19612 10896 19616
rect 10832 19556 10836 19612
rect 10836 19556 10892 19612
rect 10892 19556 10896 19612
rect 10832 19552 10896 19556
rect 10912 19612 10976 19616
rect 10912 19556 10916 19612
rect 10916 19556 10972 19612
rect 10972 19556 10976 19612
rect 10912 19552 10976 19556
rect 10992 19612 11056 19616
rect 10992 19556 10996 19612
rect 10996 19556 11052 19612
rect 11052 19556 11056 19612
rect 10992 19552 11056 19556
rect 13752 19612 13816 19616
rect 13752 19556 13756 19612
rect 13756 19556 13812 19612
rect 13812 19556 13816 19612
rect 13752 19552 13816 19556
rect 13832 19612 13896 19616
rect 13832 19556 13836 19612
rect 13836 19556 13892 19612
rect 13892 19556 13896 19612
rect 13832 19552 13896 19556
rect 13912 19612 13976 19616
rect 13912 19556 13916 19612
rect 13916 19556 13972 19612
rect 13972 19556 13976 19612
rect 13912 19552 13976 19556
rect 13992 19612 14056 19616
rect 13992 19556 13996 19612
rect 13996 19556 14052 19612
rect 14052 19556 14056 19612
rect 13992 19552 14056 19556
rect 16752 19612 16816 19616
rect 16752 19556 16756 19612
rect 16756 19556 16812 19612
rect 16812 19556 16816 19612
rect 16752 19552 16816 19556
rect 16832 19612 16896 19616
rect 16832 19556 16836 19612
rect 16836 19556 16892 19612
rect 16892 19556 16896 19612
rect 16832 19552 16896 19556
rect 16912 19612 16976 19616
rect 16912 19556 16916 19612
rect 16916 19556 16972 19612
rect 16972 19556 16976 19612
rect 16912 19552 16976 19556
rect 16992 19612 17056 19616
rect 16992 19556 16996 19612
rect 16996 19556 17052 19612
rect 17052 19556 17056 19612
rect 16992 19552 17056 19556
rect 19752 19612 19816 19616
rect 19752 19556 19756 19612
rect 19756 19556 19812 19612
rect 19812 19556 19816 19612
rect 19752 19552 19816 19556
rect 19832 19612 19896 19616
rect 19832 19556 19836 19612
rect 19836 19556 19892 19612
rect 19892 19556 19896 19612
rect 19832 19552 19896 19556
rect 19912 19612 19976 19616
rect 19912 19556 19916 19612
rect 19916 19556 19972 19612
rect 19972 19556 19976 19612
rect 19912 19552 19976 19556
rect 19992 19612 20056 19616
rect 19992 19556 19996 19612
rect 19996 19556 20052 19612
rect 20052 19556 20056 19612
rect 19992 19552 20056 19556
rect 22752 19612 22816 19616
rect 22752 19556 22756 19612
rect 22756 19556 22812 19612
rect 22812 19556 22816 19612
rect 22752 19552 22816 19556
rect 22832 19612 22896 19616
rect 22832 19556 22836 19612
rect 22836 19556 22892 19612
rect 22892 19556 22896 19612
rect 22832 19552 22896 19556
rect 22912 19612 22976 19616
rect 22912 19556 22916 19612
rect 22916 19556 22972 19612
rect 22972 19556 22976 19612
rect 22912 19552 22976 19556
rect 22992 19612 23056 19616
rect 22992 19556 22996 19612
rect 22996 19556 23052 19612
rect 23052 19556 23056 19612
rect 22992 19552 23056 19556
rect 25752 19612 25816 19616
rect 25752 19556 25756 19612
rect 25756 19556 25812 19612
rect 25812 19556 25816 19612
rect 25752 19552 25816 19556
rect 25832 19612 25896 19616
rect 25832 19556 25836 19612
rect 25836 19556 25892 19612
rect 25892 19556 25896 19612
rect 25832 19552 25896 19556
rect 25912 19612 25976 19616
rect 25912 19556 25916 19612
rect 25916 19556 25972 19612
rect 25972 19556 25976 19612
rect 25912 19552 25976 19556
rect 25992 19612 26056 19616
rect 25992 19556 25996 19612
rect 25996 19556 26052 19612
rect 26052 19556 26056 19612
rect 25992 19552 26056 19556
rect 3252 19068 3316 19072
rect 3252 19012 3256 19068
rect 3256 19012 3312 19068
rect 3312 19012 3316 19068
rect 3252 19008 3316 19012
rect 3332 19068 3396 19072
rect 3332 19012 3336 19068
rect 3336 19012 3392 19068
rect 3392 19012 3396 19068
rect 3332 19008 3396 19012
rect 3412 19068 3476 19072
rect 3412 19012 3416 19068
rect 3416 19012 3472 19068
rect 3472 19012 3476 19068
rect 3412 19008 3476 19012
rect 3492 19068 3556 19072
rect 3492 19012 3496 19068
rect 3496 19012 3552 19068
rect 3552 19012 3556 19068
rect 3492 19008 3556 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 6412 19068 6476 19072
rect 6412 19012 6416 19068
rect 6416 19012 6472 19068
rect 6472 19012 6476 19068
rect 6412 19008 6476 19012
rect 6492 19068 6556 19072
rect 6492 19012 6496 19068
rect 6496 19012 6552 19068
rect 6552 19012 6556 19068
rect 6492 19008 6556 19012
rect 9252 19068 9316 19072
rect 9252 19012 9256 19068
rect 9256 19012 9312 19068
rect 9312 19012 9316 19068
rect 9252 19008 9316 19012
rect 9332 19068 9396 19072
rect 9332 19012 9336 19068
rect 9336 19012 9392 19068
rect 9392 19012 9396 19068
rect 9332 19008 9396 19012
rect 9412 19068 9476 19072
rect 9412 19012 9416 19068
rect 9416 19012 9472 19068
rect 9472 19012 9476 19068
rect 9412 19008 9476 19012
rect 9492 19068 9556 19072
rect 9492 19012 9496 19068
rect 9496 19012 9552 19068
rect 9552 19012 9556 19068
rect 9492 19008 9556 19012
rect 12252 19068 12316 19072
rect 12252 19012 12256 19068
rect 12256 19012 12312 19068
rect 12312 19012 12316 19068
rect 12252 19008 12316 19012
rect 12332 19068 12396 19072
rect 12332 19012 12336 19068
rect 12336 19012 12392 19068
rect 12392 19012 12396 19068
rect 12332 19008 12396 19012
rect 12412 19068 12476 19072
rect 12412 19012 12416 19068
rect 12416 19012 12472 19068
rect 12472 19012 12476 19068
rect 12412 19008 12476 19012
rect 12492 19068 12556 19072
rect 12492 19012 12496 19068
rect 12496 19012 12552 19068
rect 12552 19012 12556 19068
rect 12492 19008 12556 19012
rect 15252 19068 15316 19072
rect 15252 19012 15256 19068
rect 15256 19012 15312 19068
rect 15312 19012 15316 19068
rect 15252 19008 15316 19012
rect 15332 19068 15396 19072
rect 15332 19012 15336 19068
rect 15336 19012 15392 19068
rect 15392 19012 15396 19068
rect 15332 19008 15396 19012
rect 15412 19068 15476 19072
rect 15412 19012 15416 19068
rect 15416 19012 15472 19068
rect 15472 19012 15476 19068
rect 15412 19008 15476 19012
rect 15492 19068 15556 19072
rect 15492 19012 15496 19068
rect 15496 19012 15552 19068
rect 15552 19012 15556 19068
rect 15492 19008 15556 19012
rect 18252 19068 18316 19072
rect 18252 19012 18256 19068
rect 18256 19012 18312 19068
rect 18312 19012 18316 19068
rect 18252 19008 18316 19012
rect 18332 19068 18396 19072
rect 18332 19012 18336 19068
rect 18336 19012 18392 19068
rect 18392 19012 18396 19068
rect 18332 19008 18396 19012
rect 18412 19068 18476 19072
rect 18412 19012 18416 19068
rect 18416 19012 18472 19068
rect 18472 19012 18476 19068
rect 18412 19008 18476 19012
rect 18492 19068 18556 19072
rect 18492 19012 18496 19068
rect 18496 19012 18552 19068
rect 18552 19012 18556 19068
rect 18492 19008 18556 19012
rect 21252 19068 21316 19072
rect 21252 19012 21256 19068
rect 21256 19012 21312 19068
rect 21312 19012 21316 19068
rect 21252 19008 21316 19012
rect 21332 19068 21396 19072
rect 21332 19012 21336 19068
rect 21336 19012 21392 19068
rect 21392 19012 21396 19068
rect 21332 19008 21396 19012
rect 21412 19068 21476 19072
rect 21412 19012 21416 19068
rect 21416 19012 21472 19068
rect 21472 19012 21476 19068
rect 21412 19008 21476 19012
rect 21492 19068 21556 19072
rect 21492 19012 21496 19068
rect 21496 19012 21552 19068
rect 21552 19012 21556 19068
rect 21492 19008 21556 19012
rect 24252 19068 24316 19072
rect 24252 19012 24256 19068
rect 24256 19012 24312 19068
rect 24312 19012 24316 19068
rect 24252 19008 24316 19012
rect 24332 19068 24396 19072
rect 24332 19012 24336 19068
rect 24336 19012 24392 19068
rect 24392 19012 24396 19068
rect 24332 19008 24396 19012
rect 24412 19068 24476 19072
rect 24412 19012 24416 19068
rect 24416 19012 24472 19068
rect 24472 19012 24476 19068
rect 24412 19008 24476 19012
rect 24492 19068 24556 19072
rect 24492 19012 24496 19068
rect 24496 19012 24552 19068
rect 24552 19012 24556 19068
rect 24492 19008 24556 19012
rect 27252 19068 27316 19072
rect 27252 19012 27256 19068
rect 27256 19012 27312 19068
rect 27312 19012 27316 19068
rect 27252 19008 27316 19012
rect 27332 19068 27396 19072
rect 27332 19012 27336 19068
rect 27336 19012 27392 19068
rect 27392 19012 27396 19068
rect 27332 19008 27396 19012
rect 27412 19068 27476 19072
rect 27412 19012 27416 19068
rect 27416 19012 27472 19068
rect 27472 19012 27476 19068
rect 27412 19008 27476 19012
rect 27492 19068 27556 19072
rect 27492 19012 27496 19068
rect 27496 19012 27552 19068
rect 27552 19012 27556 19068
rect 27492 19008 27556 19012
rect 1752 18524 1816 18528
rect 1752 18468 1756 18524
rect 1756 18468 1812 18524
rect 1812 18468 1816 18524
rect 1752 18464 1816 18468
rect 1832 18524 1896 18528
rect 1832 18468 1836 18524
rect 1836 18468 1892 18524
rect 1892 18468 1896 18524
rect 1832 18464 1896 18468
rect 1912 18524 1976 18528
rect 1912 18468 1916 18524
rect 1916 18468 1972 18524
rect 1972 18468 1976 18524
rect 1912 18464 1976 18468
rect 1992 18524 2056 18528
rect 1992 18468 1996 18524
rect 1996 18468 2052 18524
rect 2052 18468 2056 18524
rect 1992 18464 2056 18468
rect 4752 18524 4816 18528
rect 4752 18468 4756 18524
rect 4756 18468 4812 18524
rect 4812 18468 4816 18524
rect 4752 18464 4816 18468
rect 4832 18524 4896 18528
rect 4832 18468 4836 18524
rect 4836 18468 4892 18524
rect 4892 18468 4896 18524
rect 4832 18464 4896 18468
rect 4912 18524 4976 18528
rect 4912 18468 4916 18524
rect 4916 18468 4972 18524
rect 4972 18468 4976 18524
rect 4912 18464 4976 18468
rect 4992 18524 5056 18528
rect 4992 18468 4996 18524
rect 4996 18468 5052 18524
rect 5052 18468 5056 18524
rect 4992 18464 5056 18468
rect 7752 18524 7816 18528
rect 7752 18468 7756 18524
rect 7756 18468 7812 18524
rect 7812 18468 7816 18524
rect 7752 18464 7816 18468
rect 7832 18524 7896 18528
rect 7832 18468 7836 18524
rect 7836 18468 7892 18524
rect 7892 18468 7896 18524
rect 7832 18464 7896 18468
rect 7912 18524 7976 18528
rect 7912 18468 7916 18524
rect 7916 18468 7972 18524
rect 7972 18468 7976 18524
rect 7912 18464 7976 18468
rect 7992 18524 8056 18528
rect 7992 18468 7996 18524
rect 7996 18468 8052 18524
rect 8052 18468 8056 18524
rect 7992 18464 8056 18468
rect 10752 18524 10816 18528
rect 10752 18468 10756 18524
rect 10756 18468 10812 18524
rect 10812 18468 10816 18524
rect 10752 18464 10816 18468
rect 10832 18524 10896 18528
rect 10832 18468 10836 18524
rect 10836 18468 10892 18524
rect 10892 18468 10896 18524
rect 10832 18464 10896 18468
rect 10912 18524 10976 18528
rect 10912 18468 10916 18524
rect 10916 18468 10972 18524
rect 10972 18468 10976 18524
rect 10912 18464 10976 18468
rect 10992 18524 11056 18528
rect 10992 18468 10996 18524
rect 10996 18468 11052 18524
rect 11052 18468 11056 18524
rect 10992 18464 11056 18468
rect 13752 18524 13816 18528
rect 13752 18468 13756 18524
rect 13756 18468 13812 18524
rect 13812 18468 13816 18524
rect 13752 18464 13816 18468
rect 13832 18524 13896 18528
rect 13832 18468 13836 18524
rect 13836 18468 13892 18524
rect 13892 18468 13896 18524
rect 13832 18464 13896 18468
rect 13912 18524 13976 18528
rect 13912 18468 13916 18524
rect 13916 18468 13972 18524
rect 13972 18468 13976 18524
rect 13912 18464 13976 18468
rect 13992 18524 14056 18528
rect 13992 18468 13996 18524
rect 13996 18468 14052 18524
rect 14052 18468 14056 18524
rect 13992 18464 14056 18468
rect 16752 18524 16816 18528
rect 16752 18468 16756 18524
rect 16756 18468 16812 18524
rect 16812 18468 16816 18524
rect 16752 18464 16816 18468
rect 16832 18524 16896 18528
rect 16832 18468 16836 18524
rect 16836 18468 16892 18524
rect 16892 18468 16896 18524
rect 16832 18464 16896 18468
rect 16912 18524 16976 18528
rect 16912 18468 16916 18524
rect 16916 18468 16972 18524
rect 16972 18468 16976 18524
rect 16912 18464 16976 18468
rect 16992 18524 17056 18528
rect 16992 18468 16996 18524
rect 16996 18468 17052 18524
rect 17052 18468 17056 18524
rect 16992 18464 17056 18468
rect 19752 18524 19816 18528
rect 19752 18468 19756 18524
rect 19756 18468 19812 18524
rect 19812 18468 19816 18524
rect 19752 18464 19816 18468
rect 19832 18524 19896 18528
rect 19832 18468 19836 18524
rect 19836 18468 19892 18524
rect 19892 18468 19896 18524
rect 19832 18464 19896 18468
rect 19912 18524 19976 18528
rect 19912 18468 19916 18524
rect 19916 18468 19972 18524
rect 19972 18468 19976 18524
rect 19912 18464 19976 18468
rect 19992 18524 20056 18528
rect 19992 18468 19996 18524
rect 19996 18468 20052 18524
rect 20052 18468 20056 18524
rect 19992 18464 20056 18468
rect 22752 18524 22816 18528
rect 22752 18468 22756 18524
rect 22756 18468 22812 18524
rect 22812 18468 22816 18524
rect 22752 18464 22816 18468
rect 22832 18524 22896 18528
rect 22832 18468 22836 18524
rect 22836 18468 22892 18524
rect 22892 18468 22896 18524
rect 22832 18464 22896 18468
rect 22912 18524 22976 18528
rect 22912 18468 22916 18524
rect 22916 18468 22972 18524
rect 22972 18468 22976 18524
rect 22912 18464 22976 18468
rect 22992 18524 23056 18528
rect 22992 18468 22996 18524
rect 22996 18468 23052 18524
rect 23052 18468 23056 18524
rect 22992 18464 23056 18468
rect 25752 18524 25816 18528
rect 25752 18468 25756 18524
rect 25756 18468 25812 18524
rect 25812 18468 25816 18524
rect 25752 18464 25816 18468
rect 25832 18524 25896 18528
rect 25832 18468 25836 18524
rect 25836 18468 25892 18524
rect 25892 18468 25896 18524
rect 25832 18464 25896 18468
rect 25912 18524 25976 18528
rect 25912 18468 25916 18524
rect 25916 18468 25972 18524
rect 25972 18468 25976 18524
rect 25912 18464 25976 18468
rect 25992 18524 26056 18528
rect 25992 18468 25996 18524
rect 25996 18468 26052 18524
rect 26052 18468 26056 18524
rect 25992 18464 26056 18468
rect 3252 17980 3316 17984
rect 3252 17924 3256 17980
rect 3256 17924 3312 17980
rect 3312 17924 3316 17980
rect 3252 17920 3316 17924
rect 3332 17980 3396 17984
rect 3332 17924 3336 17980
rect 3336 17924 3392 17980
rect 3392 17924 3396 17980
rect 3332 17920 3396 17924
rect 3412 17980 3476 17984
rect 3412 17924 3416 17980
rect 3416 17924 3472 17980
rect 3472 17924 3476 17980
rect 3412 17920 3476 17924
rect 3492 17980 3556 17984
rect 3492 17924 3496 17980
rect 3496 17924 3552 17980
rect 3552 17924 3556 17980
rect 3492 17920 3556 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 6412 17980 6476 17984
rect 6412 17924 6416 17980
rect 6416 17924 6472 17980
rect 6472 17924 6476 17980
rect 6412 17920 6476 17924
rect 6492 17980 6556 17984
rect 6492 17924 6496 17980
rect 6496 17924 6552 17980
rect 6552 17924 6556 17980
rect 6492 17920 6556 17924
rect 9252 17980 9316 17984
rect 9252 17924 9256 17980
rect 9256 17924 9312 17980
rect 9312 17924 9316 17980
rect 9252 17920 9316 17924
rect 9332 17980 9396 17984
rect 9332 17924 9336 17980
rect 9336 17924 9392 17980
rect 9392 17924 9396 17980
rect 9332 17920 9396 17924
rect 9412 17980 9476 17984
rect 9412 17924 9416 17980
rect 9416 17924 9472 17980
rect 9472 17924 9476 17980
rect 9412 17920 9476 17924
rect 9492 17980 9556 17984
rect 9492 17924 9496 17980
rect 9496 17924 9552 17980
rect 9552 17924 9556 17980
rect 9492 17920 9556 17924
rect 12252 17980 12316 17984
rect 12252 17924 12256 17980
rect 12256 17924 12312 17980
rect 12312 17924 12316 17980
rect 12252 17920 12316 17924
rect 12332 17980 12396 17984
rect 12332 17924 12336 17980
rect 12336 17924 12392 17980
rect 12392 17924 12396 17980
rect 12332 17920 12396 17924
rect 12412 17980 12476 17984
rect 12412 17924 12416 17980
rect 12416 17924 12472 17980
rect 12472 17924 12476 17980
rect 12412 17920 12476 17924
rect 12492 17980 12556 17984
rect 12492 17924 12496 17980
rect 12496 17924 12552 17980
rect 12552 17924 12556 17980
rect 12492 17920 12556 17924
rect 15252 17980 15316 17984
rect 15252 17924 15256 17980
rect 15256 17924 15312 17980
rect 15312 17924 15316 17980
rect 15252 17920 15316 17924
rect 15332 17980 15396 17984
rect 15332 17924 15336 17980
rect 15336 17924 15392 17980
rect 15392 17924 15396 17980
rect 15332 17920 15396 17924
rect 15412 17980 15476 17984
rect 15412 17924 15416 17980
rect 15416 17924 15472 17980
rect 15472 17924 15476 17980
rect 15412 17920 15476 17924
rect 15492 17980 15556 17984
rect 15492 17924 15496 17980
rect 15496 17924 15552 17980
rect 15552 17924 15556 17980
rect 15492 17920 15556 17924
rect 18252 17980 18316 17984
rect 18252 17924 18256 17980
rect 18256 17924 18312 17980
rect 18312 17924 18316 17980
rect 18252 17920 18316 17924
rect 18332 17980 18396 17984
rect 18332 17924 18336 17980
rect 18336 17924 18392 17980
rect 18392 17924 18396 17980
rect 18332 17920 18396 17924
rect 18412 17980 18476 17984
rect 18412 17924 18416 17980
rect 18416 17924 18472 17980
rect 18472 17924 18476 17980
rect 18412 17920 18476 17924
rect 18492 17980 18556 17984
rect 18492 17924 18496 17980
rect 18496 17924 18552 17980
rect 18552 17924 18556 17980
rect 18492 17920 18556 17924
rect 21252 17980 21316 17984
rect 21252 17924 21256 17980
rect 21256 17924 21312 17980
rect 21312 17924 21316 17980
rect 21252 17920 21316 17924
rect 21332 17980 21396 17984
rect 21332 17924 21336 17980
rect 21336 17924 21392 17980
rect 21392 17924 21396 17980
rect 21332 17920 21396 17924
rect 21412 17980 21476 17984
rect 21412 17924 21416 17980
rect 21416 17924 21472 17980
rect 21472 17924 21476 17980
rect 21412 17920 21476 17924
rect 21492 17980 21556 17984
rect 21492 17924 21496 17980
rect 21496 17924 21552 17980
rect 21552 17924 21556 17980
rect 21492 17920 21556 17924
rect 24252 17980 24316 17984
rect 24252 17924 24256 17980
rect 24256 17924 24312 17980
rect 24312 17924 24316 17980
rect 24252 17920 24316 17924
rect 24332 17980 24396 17984
rect 24332 17924 24336 17980
rect 24336 17924 24392 17980
rect 24392 17924 24396 17980
rect 24332 17920 24396 17924
rect 24412 17980 24476 17984
rect 24412 17924 24416 17980
rect 24416 17924 24472 17980
rect 24472 17924 24476 17980
rect 24412 17920 24476 17924
rect 24492 17980 24556 17984
rect 24492 17924 24496 17980
rect 24496 17924 24552 17980
rect 24552 17924 24556 17980
rect 24492 17920 24556 17924
rect 27252 17980 27316 17984
rect 27252 17924 27256 17980
rect 27256 17924 27312 17980
rect 27312 17924 27316 17980
rect 27252 17920 27316 17924
rect 27332 17980 27396 17984
rect 27332 17924 27336 17980
rect 27336 17924 27392 17980
rect 27392 17924 27396 17980
rect 27332 17920 27396 17924
rect 27412 17980 27476 17984
rect 27412 17924 27416 17980
rect 27416 17924 27472 17980
rect 27472 17924 27476 17980
rect 27412 17920 27476 17924
rect 27492 17980 27556 17984
rect 27492 17924 27496 17980
rect 27496 17924 27552 17980
rect 27552 17924 27556 17980
rect 27492 17920 27556 17924
rect 1752 17436 1816 17440
rect 1752 17380 1756 17436
rect 1756 17380 1812 17436
rect 1812 17380 1816 17436
rect 1752 17376 1816 17380
rect 1832 17436 1896 17440
rect 1832 17380 1836 17436
rect 1836 17380 1892 17436
rect 1892 17380 1896 17436
rect 1832 17376 1896 17380
rect 1912 17436 1976 17440
rect 1912 17380 1916 17436
rect 1916 17380 1972 17436
rect 1972 17380 1976 17436
rect 1912 17376 1976 17380
rect 1992 17436 2056 17440
rect 1992 17380 1996 17436
rect 1996 17380 2052 17436
rect 2052 17380 2056 17436
rect 1992 17376 2056 17380
rect 4752 17436 4816 17440
rect 4752 17380 4756 17436
rect 4756 17380 4812 17436
rect 4812 17380 4816 17436
rect 4752 17376 4816 17380
rect 4832 17436 4896 17440
rect 4832 17380 4836 17436
rect 4836 17380 4892 17436
rect 4892 17380 4896 17436
rect 4832 17376 4896 17380
rect 4912 17436 4976 17440
rect 4912 17380 4916 17436
rect 4916 17380 4972 17436
rect 4972 17380 4976 17436
rect 4912 17376 4976 17380
rect 4992 17436 5056 17440
rect 4992 17380 4996 17436
rect 4996 17380 5052 17436
rect 5052 17380 5056 17436
rect 4992 17376 5056 17380
rect 7752 17436 7816 17440
rect 7752 17380 7756 17436
rect 7756 17380 7812 17436
rect 7812 17380 7816 17436
rect 7752 17376 7816 17380
rect 7832 17436 7896 17440
rect 7832 17380 7836 17436
rect 7836 17380 7892 17436
rect 7892 17380 7896 17436
rect 7832 17376 7896 17380
rect 7912 17436 7976 17440
rect 7912 17380 7916 17436
rect 7916 17380 7972 17436
rect 7972 17380 7976 17436
rect 7912 17376 7976 17380
rect 7992 17436 8056 17440
rect 7992 17380 7996 17436
rect 7996 17380 8052 17436
rect 8052 17380 8056 17436
rect 7992 17376 8056 17380
rect 10752 17436 10816 17440
rect 10752 17380 10756 17436
rect 10756 17380 10812 17436
rect 10812 17380 10816 17436
rect 10752 17376 10816 17380
rect 10832 17436 10896 17440
rect 10832 17380 10836 17436
rect 10836 17380 10892 17436
rect 10892 17380 10896 17436
rect 10832 17376 10896 17380
rect 10912 17436 10976 17440
rect 10912 17380 10916 17436
rect 10916 17380 10972 17436
rect 10972 17380 10976 17436
rect 10912 17376 10976 17380
rect 10992 17436 11056 17440
rect 10992 17380 10996 17436
rect 10996 17380 11052 17436
rect 11052 17380 11056 17436
rect 10992 17376 11056 17380
rect 13752 17436 13816 17440
rect 13752 17380 13756 17436
rect 13756 17380 13812 17436
rect 13812 17380 13816 17436
rect 13752 17376 13816 17380
rect 13832 17436 13896 17440
rect 13832 17380 13836 17436
rect 13836 17380 13892 17436
rect 13892 17380 13896 17436
rect 13832 17376 13896 17380
rect 13912 17436 13976 17440
rect 13912 17380 13916 17436
rect 13916 17380 13972 17436
rect 13972 17380 13976 17436
rect 13912 17376 13976 17380
rect 13992 17436 14056 17440
rect 13992 17380 13996 17436
rect 13996 17380 14052 17436
rect 14052 17380 14056 17436
rect 13992 17376 14056 17380
rect 16752 17436 16816 17440
rect 16752 17380 16756 17436
rect 16756 17380 16812 17436
rect 16812 17380 16816 17436
rect 16752 17376 16816 17380
rect 16832 17436 16896 17440
rect 16832 17380 16836 17436
rect 16836 17380 16892 17436
rect 16892 17380 16896 17436
rect 16832 17376 16896 17380
rect 16912 17436 16976 17440
rect 16912 17380 16916 17436
rect 16916 17380 16972 17436
rect 16972 17380 16976 17436
rect 16912 17376 16976 17380
rect 16992 17436 17056 17440
rect 16992 17380 16996 17436
rect 16996 17380 17052 17436
rect 17052 17380 17056 17436
rect 16992 17376 17056 17380
rect 19752 17436 19816 17440
rect 19752 17380 19756 17436
rect 19756 17380 19812 17436
rect 19812 17380 19816 17436
rect 19752 17376 19816 17380
rect 19832 17436 19896 17440
rect 19832 17380 19836 17436
rect 19836 17380 19892 17436
rect 19892 17380 19896 17436
rect 19832 17376 19896 17380
rect 19912 17436 19976 17440
rect 19912 17380 19916 17436
rect 19916 17380 19972 17436
rect 19972 17380 19976 17436
rect 19912 17376 19976 17380
rect 19992 17436 20056 17440
rect 19992 17380 19996 17436
rect 19996 17380 20052 17436
rect 20052 17380 20056 17436
rect 19992 17376 20056 17380
rect 22752 17436 22816 17440
rect 22752 17380 22756 17436
rect 22756 17380 22812 17436
rect 22812 17380 22816 17436
rect 22752 17376 22816 17380
rect 22832 17436 22896 17440
rect 22832 17380 22836 17436
rect 22836 17380 22892 17436
rect 22892 17380 22896 17436
rect 22832 17376 22896 17380
rect 22912 17436 22976 17440
rect 22912 17380 22916 17436
rect 22916 17380 22972 17436
rect 22972 17380 22976 17436
rect 22912 17376 22976 17380
rect 22992 17436 23056 17440
rect 22992 17380 22996 17436
rect 22996 17380 23052 17436
rect 23052 17380 23056 17436
rect 22992 17376 23056 17380
rect 25752 17436 25816 17440
rect 25752 17380 25756 17436
rect 25756 17380 25812 17436
rect 25812 17380 25816 17436
rect 25752 17376 25816 17380
rect 25832 17436 25896 17440
rect 25832 17380 25836 17436
rect 25836 17380 25892 17436
rect 25892 17380 25896 17436
rect 25832 17376 25896 17380
rect 25912 17436 25976 17440
rect 25912 17380 25916 17436
rect 25916 17380 25972 17436
rect 25972 17380 25976 17436
rect 25912 17376 25976 17380
rect 25992 17436 26056 17440
rect 25992 17380 25996 17436
rect 25996 17380 26052 17436
rect 26052 17380 26056 17436
rect 25992 17376 26056 17380
rect 3252 16892 3316 16896
rect 3252 16836 3256 16892
rect 3256 16836 3312 16892
rect 3312 16836 3316 16892
rect 3252 16832 3316 16836
rect 3332 16892 3396 16896
rect 3332 16836 3336 16892
rect 3336 16836 3392 16892
rect 3392 16836 3396 16892
rect 3332 16832 3396 16836
rect 3412 16892 3476 16896
rect 3412 16836 3416 16892
rect 3416 16836 3472 16892
rect 3472 16836 3476 16892
rect 3412 16832 3476 16836
rect 3492 16892 3556 16896
rect 3492 16836 3496 16892
rect 3496 16836 3552 16892
rect 3552 16836 3556 16892
rect 3492 16832 3556 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 6412 16892 6476 16896
rect 6412 16836 6416 16892
rect 6416 16836 6472 16892
rect 6472 16836 6476 16892
rect 6412 16832 6476 16836
rect 6492 16892 6556 16896
rect 6492 16836 6496 16892
rect 6496 16836 6552 16892
rect 6552 16836 6556 16892
rect 6492 16832 6556 16836
rect 9252 16892 9316 16896
rect 9252 16836 9256 16892
rect 9256 16836 9312 16892
rect 9312 16836 9316 16892
rect 9252 16832 9316 16836
rect 9332 16892 9396 16896
rect 9332 16836 9336 16892
rect 9336 16836 9392 16892
rect 9392 16836 9396 16892
rect 9332 16832 9396 16836
rect 9412 16892 9476 16896
rect 9412 16836 9416 16892
rect 9416 16836 9472 16892
rect 9472 16836 9476 16892
rect 9412 16832 9476 16836
rect 9492 16892 9556 16896
rect 9492 16836 9496 16892
rect 9496 16836 9552 16892
rect 9552 16836 9556 16892
rect 9492 16832 9556 16836
rect 12252 16892 12316 16896
rect 12252 16836 12256 16892
rect 12256 16836 12312 16892
rect 12312 16836 12316 16892
rect 12252 16832 12316 16836
rect 12332 16892 12396 16896
rect 12332 16836 12336 16892
rect 12336 16836 12392 16892
rect 12392 16836 12396 16892
rect 12332 16832 12396 16836
rect 12412 16892 12476 16896
rect 12412 16836 12416 16892
rect 12416 16836 12472 16892
rect 12472 16836 12476 16892
rect 12412 16832 12476 16836
rect 12492 16892 12556 16896
rect 12492 16836 12496 16892
rect 12496 16836 12552 16892
rect 12552 16836 12556 16892
rect 12492 16832 12556 16836
rect 15252 16892 15316 16896
rect 15252 16836 15256 16892
rect 15256 16836 15312 16892
rect 15312 16836 15316 16892
rect 15252 16832 15316 16836
rect 15332 16892 15396 16896
rect 15332 16836 15336 16892
rect 15336 16836 15392 16892
rect 15392 16836 15396 16892
rect 15332 16832 15396 16836
rect 15412 16892 15476 16896
rect 15412 16836 15416 16892
rect 15416 16836 15472 16892
rect 15472 16836 15476 16892
rect 15412 16832 15476 16836
rect 15492 16892 15556 16896
rect 15492 16836 15496 16892
rect 15496 16836 15552 16892
rect 15552 16836 15556 16892
rect 15492 16832 15556 16836
rect 18252 16892 18316 16896
rect 18252 16836 18256 16892
rect 18256 16836 18312 16892
rect 18312 16836 18316 16892
rect 18252 16832 18316 16836
rect 18332 16892 18396 16896
rect 18332 16836 18336 16892
rect 18336 16836 18392 16892
rect 18392 16836 18396 16892
rect 18332 16832 18396 16836
rect 18412 16892 18476 16896
rect 18412 16836 18416 16892
rect 18416 16836 18472 16892
rect 18472 16836 18476 16892
rect 18412 16832 18476 16836
rect 18492 16892 18556 16896
rect 18492 16836 18496 16892
rect 18496 16836 18552 16892
rect 18552 16836 18556 16892
rect 18492 16832 18556 16836
rect 21252 16892 21316 16896
rect 21252 16836 21256 16892
rect 21256 16836 21312 16892
rect 21312 16836 21316 16892
rect 21252 16832 21316 16836
rect 21332 16892 21396 16896
rect 21332 16836 21336 16892
rect 21336 16836 21392 16892
rect 21392 16836 21396 16892
rect 21332 16832 21396 16836
rect 21412 16892 21476 16896
rect 21412 16836 21416 16892
rect 21416 16836 21472 16892
rect 21472 16836 21476 16892
rect 21412 16832 21476 16836
rect 21492 16892 21556 16896
rect 21492 16836 21496 16892
rect 21496 16836 21552 16892
rect 21552 16836 21556 16892
rect 21492 16832 21556 16836
rect 24252 16892 24316 16896
rect 24252 16836 24256 16892
rect 24256 16836 24312 16892
rect 24312 16836 24316 16892
rect 24252 16832 24316 16836
rect 24332 16892 24396 16896
rect 24332 16836 24336 16892
rect 24336 16836 24392 16892
rect 24392 16836 24396 16892
rect 24332 16832 24396 16836
rect 24412 16892 24476 16896
rect 24412 16836 24416 16892
rect 24416 16836 24472 16892
rect 24472 16836 24476 16892
rect 24412 16832 24476 16836
rect 24492 16892 24556 16896
rect 24492 16836 24496 16892
rect 24496 16836 24552 16892
rect 24552 16836 24556 16892
rect 24492 16832 24556 16836
rect 27252 16892 27316 16896
rect 27252 16836 27256 16892
rect 27256 16836 27312 16892
rect 27312 16836 27316 16892
rect 27252 16832 27316 16836
rect 27332 16892 27396 16896
rect 27332 16836 27336 16892
rect 27336 16836 27392 16892
rect 27392 16836 27396 16892
rect 27332 16832 27396 16836
rect 27412 16892 27476 16896
rect 27412 16836 27416 16892
rect 27416 16836 27472 16892
rect 27472 16836 27476 16892
rect 27412 16832 27476 16836
rect 27492 16892 27556 16896
rect 27492 16836 27496 16892
rect 27496 16836 27552 16892
rect 27552 16836 27556 16892
rect 27492 16832 27556 16836
rect 1752 16348 1816 16352
rect 1752 16292 1756 16348
rect 1756 16292 1812 16348
rect 1812 16292 1816 16348
rect 1752 16288 1816 16292
rect 1832 16348 1896 16352
rect 1832 16292 1836 16348
rect 1836 16292 1892 16348
rect 1892 16292 1896 16348
rect 1832 16288 1896 16292
rect 1912 16348 1976 16352
rect 1912 16292 1916 16348
rect 1916 16292 1972 16348
rect 1972 16292 1976 16348
rect 1912 16288 1976 16292
rect 1992 16348 2056 16352
rect 1992 16292 1996 16348
rect 1996 16292 2052 16348
rect 2052 16292 2056 16348
rect 1992 16288 2056 16292
rect 4752 16348 4816 16352
rect 4752 16292 4756 16348
rect 4756 16292 4812 16348
rect 4812 16292 4816 16348
rect 4752 16288 4816 16292
rect 4832 16348 4896 16352
rect 4832 16292 4836 16348
rect 4836 16292 4892 16348
rect 4892 16292 4896 16348
rect 4832 16288 4896 16292
rect 4912 16348 4976 16352
rect 4912 16292 4916 16348
rect 4916 16292 4972 16348
rect 4972 16292 4976 16348
rect 4912 16288 4976 16292
rect 4992 16348 5056 16352
rect 4992 16292 4996 16348
rect 4996 16292 5052 16348
rect 5052 16292 5056 16348
rect 4992 16288 5056 16292
rect 7752 16348 7816 16352
rect 7752 16292 7756 16348
rect 7756 16292 7812 16348
rect 7812 16292 7816 16348
rect 7752 16288 7816 16292
rect 7832 16348 7896 16352
rect 7832 16292 7836 16348
rect 7836 16292 7892 16348
rect 7892 16292 7896 16348
rect 7832 16288 7896 16292
rect 7912 16348 7976 16352
rect 7912 16292 7916 16348
rect 7916 16292 7972 16348
rect 7972 16292 7976 16348
rect 7912 16288 7976 16292
rect 7992 16348 8056 16352
rect 7992 16292 7996 16348
rect 7996 16292 8052 16348
rect 8052 16292 8056 16348
rect 7992 16288 8056 16292
rect 10752 16348 10816 16352
rect 10752 16292 10756 16348
rect 10756 16292 10812 16348
rect 10812 16292 10816 16348
rect 10752 16288 10816 16292
rect 10832 16348 10896 16352
rect 10832 16292 10836 16348
rect 10836 16292 10892 16348
rect 10892 16292 10896 16348
rect 10832 16288 10896 16292
rect 10912 16348 10976 16352
rect 10912 16292 10916 16348
rect 10916 16292 10972 16348
rect 10972 16292 10976 16348
rect 10912 16288 10976 16292
rect 10992 16348 11056 16352
rect 10992 16292 10996 16348
rect 10996 16292 11052 16348
rect 11052 16292 11056 16348
rect 10992 16288 11056 16292
rect 13752 16348 13816 16352
rect 13752 16292 13756 16348
rect 13756 16292 13812 16348
rect 13812 16292 13816 16348
rect 13752 16288 13816 16292
rect 13832 16348 13896 16352
rect 13832 16292 13836 16348
rect 13836 16292 13892 16348
rect 13892 16292 13896 16348
rect 13832 16288 13896 16292
rect 13912 16348 13976 16352
rect 13912 16292 13916 16348
rect 13916 16292 13972 16348
rect 13972 16292 13976 16348
rect 13912 16288 13976 16292
rect 13992 16348 14056 16352
rect 13992 16292 13996 16348
rect 13996 16292 14052 16348
rect 14052 16292 14056 16348
rect 13992 16288 14056 16292
rect 16752 16348 16816 16352
rect 16752 16292 16756 16348
rect 16756 16292 16812 16348
rect 16812 16292 16816 16348
rect 16752 16288 16816 16292
rect 16832 16348 16896 16352
rect 16832 16292 16836 16348
rect 16836 16292 16892 16348
rect 16892 16292 16896 16348
rect 16832 16288 16896 16292
rect 16912 16348 16976 16352
rect 16912 16292 16916 16348
rect 16916 16292 16972 16348
rect 16972 16292 16976 16348
rect 16912 16288 16976 16292
rect 16992 16348 17056 16352
rect 16992 16292 16996 16348
rect 16996 16292 17052 16348
rect 17052 16292 17056 16348
rect 16992 16288 17056 16292
rect 19752 16348 19816 16352
rect 19752 16292 19756 16348
rect 19756 16292 19812 16348
rect 19812 16292 19816 16348
rect 19752 16288 19816 16292
rect 19832 16348 19896 16352
rect 19832 16292 19836 16348
rect 19836 16292 19892 16348
rect 19892 16292 19896 16348
rect 19832 16288 19896 16292
rect 19912 16348 19976 16352
rect 19912 16292 19916 16348
rect 19916 16292 19972 16348
rect 19972 16292 19976 16348
rect 19912 16288 19976 16292
rect 19992 16348 20056 16352
rect 19992 16292 19996 16348
rect 19996 16292 20052 16348
rect 20052 16292 20056 16348
rect 19992 16288 20056 16292
rect 22752 16348 22816 16352
rect 22752 16292 22756 16348
rect 22756 16292 22812 16348
rect 22812 16292 22816 16348
rect 22752 16288 22816 16292
rect 22832 16348 22896 16352
rect 22832 16292 22836 16348
rect 22836 16292 22892 16348
rect 22892 16292 22896 16348
rect 22832 16288 22896 16292
rect 22912 16348 22976 16352
rect 22912 16292 22916 16348
rect 22916 16292 22972 16348
rect 22972 16292 22976 16348
rect 22912 16288 22976 16292
rect 22992 16348 23056 16352
rect 22992 16292 22996 16348
rect 22996 16292 23052 16348
rect 23052 16292 23056 16348
rect 22992 16288 23056 16292
rect 25752 16348 25816 16352
rect 25752 16292 25756 16348
rect 25756 16292 25812 16348
rect 25812 16292 25816 16348
rect 25752 16288 25816 16292
rect 25832 16348 25896 16352
rect 25832 16292 25836 16348
rect 25836 16292 25892 16348
rect 25892 16292 25896 16348
rect 25832 16288 25896 16292
rect 25912 16348 25976 16352
rect 25912 16292 25916 16348
rect 25916 16292 25972 16348
rect 25972 16292 25976 16348
rect 25912 16288 25976 16292
rect 25992 16348 26056 16352
rect 25992 16292 25996 16348
rect 25996 16292 26052 16348
rect 26052 16292 26056 16348
rect 25992 16288 26056 16292
rect 3252 15804 3316 15808
rect 3252 15748 3256 15804
rect 3256 15748 3312 15804
rect 3312 15748 3316 15804
rect 3252 15744 3316 15748
rect 3332 15804 3396 15808
rect 3332 15748 3336 15804
rect 3336 15748 3392 15804
rect 3392 15748 3396 15804
rect 3332 15744 3396 15748
rect 3412 15804 3476 15808
rect 3412 15748 3416 15804
rect 3416 15748 3472 15804
rect 3472 15748 3476 15804
rect 3412 15744 3476 15748
rect 3492 15804 3556 15808
rect 3492 15748 3496 15804
rect 3496 15748 3552 15804
rect 3552 15748 3556 15804
rect 3492 15744 3556 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 6412 15804 6476 15808
rect 6412 15748 6416 15804
rect 6416 15748 6472 15804
rect 6472 15748 6476 15804
rect 6412 15744 6476 15748
rect 6492 15804 6556 15808
rect 6492 15748 6496 15804
rect 6496 15748 6552 15804
rect 6552 15748 6556 15804
rect 6492 15744 6556 15748
rect 9252 15804 9316 15808
rect 9252 15748 9256 15804
rect 9256 15748 9312 15804
rect 9312 15748 9316 15804
rect 9252 15744 9316 15748
rect 9332 15804 9396 15808
rect 9332 15748 9336 15804
rect 9336 15748 9392 15804
rect 9392 15748 9396 15804
rect 9332 15744 9396 15748
rect 9412 15804 9476 15808
rect 9412 15748 9416 15804
rect 9416 15748 9472 15804
rect 9472 15748 9476 15804
rect 9412 15744 9476 15748
rect 9492 15804 9556 15808
rect 9492 15748 9496 15804
rect 9496 15748 9552 15804
rect 9552 15748 9556 15804
rect 9492 15744 9556 15748
rect 12252 15804 12316 15808
rect 12252 15748 12256 15804
rect 12256 15748 12312 15804
rect 12312 15748 12316 15804
rect 12252 15744 12316 15748
rect 12332 15804 12396 15808
rect 12332 15748 12336 15804
rect 12336 15748 12392 15804
rect 12392 15748 12396 15804
rect 12332 15744 12396 15748
rect 12412 15804 12476 15808
rect 12412 15748 12416 15804
rect 12416 15748 12472 15804
rect 12472 15748 12476 15804
rect 12412 15744 12476 15748
rect 12492 15804 12556 15808
rect 12492 15748 12496 15804
rect 12496 15748 12552 15804
rect 12552 15748 12556 15804
rect 12492 15744 12556 15748
rect 15252 15804 15316 15808
rect 15252 15748 15256 15804
rect 15256 15748 15312 15804
rect 15312 15748 15316 15804
rect 15252 15744 15316 15748
rect 15332 15804 15396 15808
rect 15332 15748 15336 15804
rect 15336 15748 15392 15804
rect 15392 15748 15396 15804
rect 15332 15744 15396 15748
rect 15412 15804 15476 15808
rect 15412 15748 15416 15804
rect 15416 15748 15472 15804
rect 15472 15748 15476 15804
rect 15412 15744 15476 15748
rect 15492 15804 15556 15808
rect 15492 15748 15496 15804
rect 15496 15748 15552 15804
rect 15552 15748 15556 15804
rect 15492 15744 15556 15748
rect 18252 15804 18316 15808
rect 18252 15748 18256 15804
rect 18256 15748 18312 15804
rect 18312 15748 18316 15804
rect 18252 15744 18316 15748
rect 18332 15804 18396 15808
rect 18332 15748 18336 15804
rect 18336 15748 18392 15804
rect 18392 15748 18396 15804
rect 18332 15744 18396 15748
rect 18412 15804 18476 15808
rect 18412 15748 18416 15804
rect 18416 15748 18472 15804
rect 18472 15748 18476 15804
rect 18412 15744 18476 15748
rect 18492 15804 18556 15808
rect 18492 15748 18496 15804
rect 18496 15748 18552 15804
rect 18552 15748 18556 15804
rect 18492 15744 18556 15748
rect 21252 15804 21316 15808
rect 21252 15748 21256 15804
rect 21256 15748 21312 15804
rect 21312 15748 21316 15804
rect 21252 15744 21316 15748
rect 21332 15804 21396 15808
rect 21332 15748 21336 15804
rect 21336 15748 21392 15804
rect 21392 15748 21396 15804
rect 21332 15744 21396 15748
rect 21412 15804 21476 15808
rect 21412 15748 21416 15804
rect 21416 15748 21472 15804
rect 21472 15748 21476 15804
rect 21412 15744 21476 15748
rect 21492 15804 21556 15808
rect 21492 15748 21496 15804
rect 21496 15748 21552 15804
rect 21552 15748 21556 15804
rect 21492 15744 21556 15748
rect 24252 15804 24316 15808
rect 24252 15748 24256 15804
rect 24256 15748 24312 15804
rect 24312 15748 24316 15804
rect 24252 15744 24316 15748
rect 24332 15804 24396 15808
rect 24332 15748 24336 15804
rect 24336 15748 24392 15804
rect 24392 15748 24396 15804
rect 24332 15744 24396 15748
rect 24412 15804 24476 15808
rect 24412 15748 24416 15804
rect 24416 15748 24472 15804
rect 24472 15748 24476 15804
rect 24412 15744 24476 15748
rect 24492 15804 24556 15808
rect 24492 15748 24496 15804
rect 24496 15748 24552 15804
rect 24552 15748 24556 15804
rect 24492 15744 24556 15748
rect 27252 15804 27316 15808
rect 27252 15748 27256 15804
rect 27256 15748 27312 15804
rect 27312 15748 27316 15804
rect 27252 15744 27316 15748
rect 27332 15804 27396 15808
rect 27332 15748 27336 15804
rect 27336 15748 27392 15804
rect 27392 15748 27396 15804
rect 27332 15744 27396 15748
rect 27412 15804 27476 15808
rect 27412 15748 27416 15804
rect 27416 15748 27472 15804
rect 27472 15748 27476 15804
rect 27412 15744 27476 15748
rect 27492 15804 27556 15808
rect 27492 15748 27496 15804
rect 27496 15748 27552 15804
rect 27552 15748 27556 15804
rect 27492 15744 27556 15748
rect 1752 15260 1816 15264
rect 1752 15204 1756 15260
rect 1756 15204 1812 15260
rect 1812 15204 1816 15260
rect 1752 15200 1816 15204
rect 1832 15260 1896 15264
rect 1832 15204 1836 15260
rect 1836 15204 1892 15260
rect 1892 15204 1896 15260
rect 1832 15200 1896 15204
rect 1912 15260 1976 15264
rect 1912 15204 1916 15260
rect 1916 15204 1972 15260
rect 1972 15204 1976 15260
rect 1912 15200 1976 15204
rect 1992 15260 2056 15264
rect 1992 15204 1996 15260
rect 1996 15204 2052 15260
rect 2052 15204 2056 15260
rect 1992 15200 2056 15204
rect 4752 15260 4816 15264
rect 4752 15204 4756 15260
rect 4756 15204 4812 15260
rect 4812 15204 4816 15260
rect 4752 15200 4816 15204
rect 4832 15260 4896 15264
rect 4832 15204 4836 15260
rect 4836 15204 4892 15260
rect 4892 15204 4896 15260
rect 4832 15200 4896 15204
rect 4912 15260 4976 15264
rect 4912 15204 4916 15260
rect 4916 15204 4972 15260
rect 4972 15204 4976 15260
rect 4912 15200 4976 15204
rect 4992 15260 5056 15264
rect 4992 15204 4996 15260
rect 4996 15204 5052 15260
rect 5052 15204 5056 15260
rect 4992 15200 5056 15204
rect 7752 15260 7816 15264
rect 7752 15204 7756 15260
rect 7756 15204 7812 15260
rect 7812 15204 7816 15260
rect 7752 15200 7816 15204
rect 7832 15260 7896 15264
rect 7832 15204 7836 15260
rect 7836 15204 7892 15260
rect 7892 15204 7896 15260
rect 7832 15200 7896 15204
rect 7912 15260 7976 15264
rect 7912 15204 7916 15260
rect 7916 15204 7972 15260
rect 7972 15204 7976 15260
rect 7912 15200 7976 15204
rect 7992 15260 8056 15264
rect 7992 15204 7996 15260
rect 7996 15204 8052 15260
rect 8052 15204 8056 15260
rect 7992 15200 8056 15204
rect 10752 15260 10816 15264
rect 10752 15204 10756 15260
rect 10756 15204 10812 15260
rect 10812 15204 10816 15260
rect 10752 15200 10816 15204
rect 10832 15260 10896 15264
rect 10832 15204 10836 15260
rect 10836 15204 10892 15260
rect 10892 15204 10896 15260
rect 10832 15200 10896 15204
rect 10912 15260 10976 15264
rect 10912 15204 10916 15260
rect 10916 15204 10972 15260
rect 10972 15204 10976 15260
rect 10912 15200 10976 15204
rect 10992 15260 11056 15264
rect 10992 15204 10996 15260
rect 10996 15204 11052 15260
rect 11052 15204 11056 15260
rect 10992 15200 11056 15204
rect 13752 15260 13816 15264
rect 13752 15204 13756 15260
rect 13756 15204 13812 15260
rect 13812 15204 13816 15260
rect 13752 15200 13816 15204
rect 13832 15260 13896 15264
rect 13832 15204 13836 15260
rect 13836 15204 13892 15260
rect 13892 15204 13896 15260
rect 13832 15200 13896 15204
rect 13912 15260 13976 15264
rect 13912 15204 13916 15260
rect 13916 15204 13972 15260
rect 13972 15204 13976 15260
rect 13912 15200 13976 15204
rect 13992 15260 14056 15264
rect 13992 15204 13996 15260
rect 13996 15204 14052 15260
rect 14052 15204 14056 15260
rect 13992 15200 14056 15204
rect 16752 15260 16816 15264
rect 16752 15204 16756 15260
rect 16756 15204 16812 15260
rect 16812 15204 16816 15260
rect 16752 15200 16816 15204
rect 16832 15260 16896 15264
rect 16832 15204 16836 15260
rect 16836 15204 16892 15260
rect 16892 15204 16896 15260
rect 16832 15200 16896 15204
rect 16912 15260 16976 15264
rect 16912 15204 16916 15260
rect 16916 15204 16972 15260
rect 16972 15204 16976 15260
rect 16912 15200 16976 15204
rect 16992 15260 17056 15264
rect 16992 15204 16996 15260
rect 16996 15204 17052 15260
rect 17052 15204 17056 15260
rect 16992 15200 17056 15204
rect 19752 15260 19816 15264
rect 19752 15204 19756 15260
rect 19756 15204 19812 15260
rect 19812 15204 19816 15260
rect 19752 15200 19816 15204
rect 19832 15260 19896 15264
rect 19832 15204 19836 15260
rect 19836 15204 19892 15260
rect 19892 15204 19896 15260
rect 19832 15200 19896 15204
rect 19912 15260 19976 15264
rect 19912 15204 19916 15260
rect 19916 15204 19972 15260
rect 19972 15204 19976 15260
rect 19912 15200 19976 15204
rect 19992 15260 20056 15264
rect 19992 15204 19996 15260
rect 19996 15204 20052 15260
rect 20052 15204 20056 15260
rect 19992 15200 20056 15204
rect 22752 15260 22816 15264
rect 22752 15204 22756 15260
rect 22756 15204 22812 15260
rect 22812 15204 22816 15260
rect 22752 15200 22816 15204
rect 22832 15260 22896 15264
rect 22832 15204 22836 15260
rect 22836 15204 22892 15260
rect 22892 15204 22896 15260
rect 22832 15200 22896 15204
rect 22912 15260 22976 15264
rect 22912 15204 22916 15260
rect 22916 15204 22972 15260
rect 22972 15204 22976 15260
rect 22912 15200 22976 15204
rect 22992 15260 23056 15264
rect 22992 15204 22996 15260
rect 22996 15204 23052 15260
rect 23052 15204 23056 15260
rect 22992 15200 23056 15204
rect 25752 15260 25816 15264
rect 25752 15204 25756 15260
rect 25756 15204 25812 15260
rect 25812 15204 25816 15260
rect 25752 15200 25816 15204
rect 25832 15260 25896 15264
rect 25832 15204 25836 15260
rect 25836 15204 25892 15260
rect 25892 15204 25896 15260
rect 25832 15200 25896 15204
rect 25912 15260 25976 15264
rect 25912 15204 25916 15260
rect 25916 15204 25972 15260
rect 25972 15204 25976 15260
rect 25912 15200 25976 15204
rect 25992 15260 26056 15264
rect 25992 15204 25996 15260
rect 25996 15204 26052 15260
rect 26052 15204 26056 15260
rect 25992 15200 26056 15204
rect 3252 14716 3316 14720
rect 3252 14660 3256 14716
rect 3256 14660 3312 14716
rect 3312 14660 3316 14716
rect 3252 14656 3316 14660
rect 3332 14716 3396 14720
rect 3332 14660 3336 14716
rect 3336 14660 3392 14716
rect 3392 14660 3396 14716
rect 3332 14656 3396 14660
rect 3412 14716 3476 14720
rect 3412 14660 3416 14716
rect 3416 14660 3472 14716
rect 3472 14660 3476 14716
rect 3412 14656 3476 14660
rect 3492 14716 3556 14720
rect 3492 14660 3496 14716
rect 3496 14660 3552 14716
rect 3552 14660 3556 14716
rect 3492 14656 3556 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 6412 14716 6476 14720
rect 6412 14660 6416 14716
rect 6416 14660 6472 14716
rect 6472 14660 6476 14716
rect 6412 14656 6476 14660
rect 6492 14716 6556 14720
rect 6492 14660 6496 14716
rect 6496 14660 6552 14716
rect 6552 14660 6556 14716
rect 6492 14656 6556 14660
rect 9252 14716 9316 14720
rect 9252 14660 9256 14716
rect 9256 14660 9312 14716
rect 9312 14660 9316 14716
rect 9252 14656 9316 14660
rect 9332 14716 9396 14720
rect 9332 14660 9336 14716
rect 9336 14660 9392 14716
rect 9392 14660 9396 14716
rect 9332 14656 9396 14660
rect 9412 14716 9476 14720
rect 9412 14660 9416 14716
rect 9416 14660 9472 14716
rect 9472 14660 9476 14716
rect 9412 14656 9476 14660
rect 9492 14716 9556 14720
rect 9492 14660 9496 14716
rect 9496 14660 9552 14716
rect 9552 14660 9556 14716
rect 9492 14656 9556 14660
rect 12252 14716 12316 14720
rect 12252 14660 12256 14716
rect 12256 14660 12312 14716
rect 12312 14660 12316 14716
rect 12252 14656 12316 14660
rect 12332 14716 12396 14720
rect 12332 14660 12336 14716
rect 12336 14660 12392 14716
rect 12392 14660 12396 14716
rect 12332 14656 12396 14660
rect 12412 14716 12476 14720
rect 12412 14660 12416 14716
rect 12416 14660 12472 14716
rect 12472 14660 12476 14716
rect 12412 14656 12476 14660
rect 12492 14716 12556 14720
rect 12492 14660 12496 14716
rect 12496 14660 12552 14716
rect 12552 14660 12556 14716
rect 12492 14656 12556 14660
rect 15252 14716 15316 14720
rect 15252 14660 15256 14716
rect 15256 14660 15312 14716
rect 15312 14660 15316 14716
rect 15252 14656 15316 14660
rect 15332 14716 15396 14720
rect 15332 14660 15336 14716
rect 15336 14660 15392 14716
rect 15392 14660 15396 14716
rect 15332 14656 15396 14660
rect 15412 14716 15476 14720
rect 15412 14660 15416 14716
rect 15416 14660 15472 14716
rect 15472 14660 15476 14716
rect 15412 14656 15476 14660
rect 15492 14716 15556 14720
rect 15492 14660 15496 14716
rect 15496 14660 15552 14716
rect 15552 14660 15556 14716
rect 15492 14656 15556 14660
rect 18252 14716 18316 14720
rect 18252 14660 18256 14716
rect 18256 14660 18312 14716
rect 18312 14660 18316 14716
rect 18252 14656 18316 14660
rect 18332 14716 18396 14720
rect 18332 14660 18336 14716
rect 18336 14660 18392 14716
rect 18392 14660 18396 14716
rect 18332 14656 18396 14660
rect 18412 14716 18476 14720
rect 18412 14660 18416 14716
rect 18416 14660 18472 14716
rect 18472 14660 18476 14716
rect 18412 14656 18476 14660
rect 18492 14716 18556 14720
rect 18492 14660 18496 14716
rect 18496 14660 18552 14716
rect 18552 14660 18556 14716
rect 18492 14656 18556 14660
rect 21252 14716 21316 14720
rect 21252 14660 21256 14716
rect 21256 14660 21312 14716
rect 21312 14660 21316 14716
rect 21252 14656 21316 14660
rect 21332 14716 21396 14720
rect 21332 14660 21336 14716
rect 21336 14660 21392 14716
rect 21392 14660 21396 14716
rect 21332 14656 21396 14660
rect 21412 14716 21476 14720
rect 21412 14660 21416 14716
rect 21416 14660 21472 14716
rect 21472 14660 21476 14716
rect 21412 14656 21476 14660
rect 21492 14716 21556 14720
rect 21492 14660 21496 14716
rect 21496 14660 21552 14716
rect 21552 14660 21556 14716
rect 21492 14656 21556 14660
rect 24252 14716 24316 14720
rect 24252 14660 24256 14716
rect 24256 14660 24312 14716
rect 24312 14660 24316 14716
rect 24252 14656 24316 14660
rect 24332 14716 24396 14720
rect 24332 14660 24336 14716
rect 24336 14660 24392 14716
rect 24392 14660 24396 14716
rect 24332 14656 24396 14660
rect 24412 14716 24476 14720
rect 24412 14660 24416 14716
rect 24416 14660 24472 14716
rect 24472 14660 24476 14716
rect 24412 14656 24476 14660
rect 24492 14716 24556 14720
rect 24492 14660 24496 14716
rect 24496 14660 24552 14716
rect 24552 14660 24556 14716
rect 24492 14656 24556 14660
rect 27252 14716 27316 14720
rect 27252 14660 27256 14716
rect 27256 14660 27312 14716
rect 27312 14660 27316 14716
rect 27252 14656 27316 14660
rect 27332 14716 27396 14720
rect 27332 14660 27336 14716
rect 27336 14660 27392 14716
rect 27392 14660 27396 14716
rect 27332 14656 27396 14660
rect 27412 14716 27476 14720
rect 27412 14660 27416 14716
rect 27416 14660 27472 14716
rect 27472 14660 27476 14716
rect 27412 14656 27476 14660
rect 27492 14716 27556 14720
rect 27492 14660 27496 14716
rect 27496 14660 27552 14716
rect 27552 14660 27556 14716
rect 27492 14656 27556 14660
rect 19380 14452 19444 14516
rect 1752 14172 1816 14176
rect 1752 14116 1756 14172
rect 1756 14116 1812 14172
rect 1812 14116 1816 14172
rect 1752 14112 1816 14116
rect 1832 14172 1896 14176
rect 1832 14116 1836 14172
rect 1836 14116 1892 14172
rect 1892 14116 1896 14172
rect 1832 14112 1896 14116
rect 1912 14172 1976 14176
rect 1912 14116 1916 14172
rect 1916 14116 1972 14172
rect 1972 14116 1976 14172
rect 1912 14112 1976 14116
rect 1992 14172 2056 14176
rect 1992 14116 1996 14172
rect 1996 14116 2052 14172
rect 2052 14116 2056 14172
rect 1992 14112 2056 14116
rect 4752 14172 4816 14176
rect 4752 14116 4756 14172
rect 4756 14116 4812 14172
rect 4812 14116 4816 14172
rect 4752 14112 4816 14116
rect 4832 14172 4896 14176
rect 4832 14116 4836 14172
rect 4836 14116 4892 14172
rect 4892 14116 4896 14172
rect 4832 14112 4896 14116
rect 4912 14172 4976 14176
rect 4912 14116 4916 14172
rect 4916 14116 4972 14172
rect 4972 14116 4976 14172
rect 4912 14112 4976 14116
rect 4992 14172 5056 14176
rect 4992 14116 4996 14172
rect 4996 14116 5052 14172
rect 5052 14116 5056 14172
rect 4992 14112 5056 14116
rect 7752 14172 7816 14176
rect 7752 14116 7756 14172
rect 7756 14116 7812 14172
rect 7812 14116 7816 14172
rect 7752 14112 7816 14116
rect 7832 14172 7896 14176
rect 7832 14116 7836 14172
rect 7836 14116 7892 14172
rect 7892 14116 7896 14172
rect 7832 14112 7896 14116
rect 7912 14172 7976 14176
rect 7912 14116 7916 14172
rect 7916 14116 7972 14172
rect 7972 14116 7976 14172
rect 7912 14112 7976 14116
rect 7992 14172 8056 14176
rect 7992 14116 7996 14172
rect 7996 14116 8052 14172
rect 8052 14116 8056 14172
rect 7992 14112 8056 14116
rect 10752 14172 10816 14176
rect 10752 14116 10756 14172
rect 10756 14116 10812 14172
rect 10812 14116 10816 14172
rect 10752 14112 10816 14116
rect 10832 14172 10896 14176
rect 10832 14116 10836 14172
rect 10836 14116 10892 14172
rect 10892 14116 10896 14172
rect 10832 14112 10896 14116
rect 10912 14172 10976 14176
rect 10912 14116 10916 14172
rect 10916 14116 10972 14172
rect 10972 14116 10976 14172
rect 10912 14112 10976 14116
rect 10992 14172 11056 14176
rect 10992 14116 10996 14172
rect 10996 14116 11052 14172
rect 11052 14116 11056 14172
rect 10992 14112 11056 14116
rect 13752 14172 13816 14176
rect 13752 14116 13756 14172
rect 13756 14116 13812 14172
rect 13812 14116 13816 14172
rect 13752 14112 13816 14116
rect 13832 14172 13896 14176
rect 13832 14116 13836 14172
rect 13836 14116 13892 14172
rect 13892 14116 13896 14172
rect 13832 14112 13896 14116
rect 13912 14172 13976 14176
rect 13912 14116 13916 14172
rect 13916 14116 13972 14172
rect 13972 14116 13976 14172
rect 13912 14112 13976 14116
rect 13992 14172 14056 14176
rect 13992 14116 13996 14172
rect 13996 14116 14052 14172
rect 14052 14116 14056 14172
rect 13992 14112 14056 14116
rect 16752 14172 16816 14176
rect 16752 14116 16756 14172
rect 16756 14116 16812 14172
rect 16812 14116 16816 14172
rect 16752 14112 16816 14116
rect 16832 14172 16896 14176
rect 16832 14116 16836 14172
rect 16836 14116 16892 14172
rect 16892 14116 16896 14172
rect 16832 14112 16896 14116
rect 16912 14172 16976 14176
rect 16912 14116 16916 14172
rect 16916 14116 16972 14172
rect 16972 14116 16976 14172
rect 16912 14112 16976 14116
rect 16992 14172 17056 14176
rect 16992 14116 16996 14172
rect 16996 14116 17052 14172
rect 17052 14116 17056 14172
rect 16992 14112 17056 14116
rect 19752 14172 19816 14176
rect 19752 14116 19756 14172
rect 19756 14116 19812 14172
rect 19812 14116 19816 14172
rect 19752 14112 19816 14116
rect 19832 14172 19896 14176
rect 19832 14116 19836 14172
rect 19836 14116 19892 14172
rect 19892 14116 19896 14172
rect 19832 14112 19896 14116
rect 19912 14172 19976 14176
rect 19912 14116 19916 14172
rect 19916 14116 19972 14172
rect 19972 14116 19976 14172
rect 19912 14112 19976 14116
rect 19992 14172 20056 14176
rect 19992 14116 19996 14172
rect 19996 14116 20052 14172
rect 20052 14116 20056 14172
rect 19992 14112 20056 14116
rect 22752 14172 22816 14176
rect 22752 14116 22756 14172
rect 22756 14116 22812 14172
rect 22812 14116 22816 14172
rect 22752 14112 22816 14116
rect 22832 14172 22896 14176
rect 22832 14116 22836 14172
rect 22836 14116 22892 14172
rect 22892 14116 22896 14172
rect 22832 14112 22896 14116
rect 22912 14172 22976 14176
rect 22912 14116 22916 14172
rect 22916 14116 22972 14172
rect 22972 14116 22976 14172
rect 22912 14112 22976 14116
rect 22992 14172 23056 14176
rect 22992 14116 22996 14172
rect 22996 14116 23052 14172
rect 23052 14116 23056 14172
rect 22992 14112 23056 14116
rect 25752 14172 25816 14176
rect 25752 14116 25756 14172
rect 25756 14116 25812 14172
rect 25812 14116 25816 14172
rect 25752 14112 25816 14116
rect 25832 14172 25896 14176
rect 25832 14116 25836 14172
rect 25836 14116 25892 14172
rect 25892 14116 25896 14172
rect 25832 14112 25896 14116
rect 25912 14172 25976 14176
rect 25912 14116 25916 14172
rect 25916 14116 25972 14172
rect 25972 14116 25976 14172
rect 25912 14112 25976 14116
rect 25992 14172 26056 14176
rect 25992 14116 25996 14172
rect 25996 14116 26052 14172
rect 26052 14116 26056 14172
rect 25992 14112 26056 14116
rect 3252 13628 3316 13632
rect 3252 13572 3256 13628
rect 3256 13572 3312 13628
rect 3312 13572 3316 13628
rect 3252 13568 3316 13572
rect 3332 13628 3396 13632
rect 3332 13572 3336 13628
rect 3336 13572 3392 13628
rect 3392 13572 3396 13628
rect 3332 13568 3396 13572
rect 3412 13628 3476 13632
rect 3412 13572 3416 13628
rect 3416 13572 3472 13628
rect 3472 13572 3476 13628
rect 3412 13568 3476 13572
rect 3492 13628 3556 13632
rect 3492 13572 3496 13628
rect 3496 13572 3552 13628
rect 3552 13572 3556 13628
rect 3492 13568 3556 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 6412 13628 6476 13632
rect 6412 13572 6416 13628
rect 6416 13572 6472 13628
rect 6472 13572 6476 13628
rect 6412 13568 6476 13572
rect 6492 13628 6556 13632
rect 6492 13572 6496 13628
rect 6496 13572 6552 13628
rect 6552 13572 6556 13628
rect 6492 13568 6556 13572
rect 9252 13628 9316 13632
rect 9252 13572 9256 13628
rect 9256 13572 9312 13628
rect 9312 13572 9316 13628
rect 9252 13568 9316 13572
rect 9332 13628 9396 13632
rect 9332 13572 9336 13628
rect 9336 13572 9392 13628
rect 9392 13572 9396 13628
rect 9332 13568 9396 13572
rect 9412 13628 9476 13632
rect 9412 13572 9416 13628
rect 9416 13572 9472 13628
rect 9472 13572 9476 13628
rect 9412 13568 9476 13572
rect 9492 13628 9556 13632
rect 9492 13572 9496 13628
rect 9496 13572 9552 13628
rect 9552 13572 9556 13628
rect 9492 13568 9556 13572
rect 12252 13628 12316 13632
rect 12252 13572 12256 13628
rect 12256 13572 12312 13628
rect 12312 13572 12316 13628
rect 12252 13568 12316 13572
rect 12332 13628 12396 13632
rect 12332 13572 12336 13628
rect 12336 13572 12392 13628
rect 12392 13572 12396 13628
rect 12332 13568 12396 13572
rect 12412 13628 12476 13632
rect 12412 13572 12416 13628
rect 12416 13572 12472 13628
rect 12472 13572 12476 13628
rect 12412 13568 12476 13572
rect 12492 13628 12556 13632
rect 12492 13572 12496 13628
rect 12496 13572 12552 13628
rect 12552 13572 12556 13628
rect 12492 13568 12556 13572
rect 15252 13628 15316 13632
rect 15252 13572 15256 13628
rect 15256 13572 15312 13628
rect 15312 13572 15316 13628
rect 15252 13568 15316 13572
rect 15332 13628 15396 13632
rect 15332 13572 15336 13628
rect 15336 13572 15392 13628
rect 15392 13572 15396 13628
rect 15332 13568 15396 13572
rect 15412 13628 15476 13632
rect 15412 13572 15416 13628
rect 15416 13572 15472 13628
rect 15472 13572 15476 13628
rect 15412 13568 15476 13572
rect 15492 13628 15556 13632
rect 15492 13572 15496 13628
rect 15496 13572 15552 13628
rect 15552 13572 15556 13628
rect 15492 13568 15556 13572
rect 18252 13628 18316 13632
rect 18252 13572 18256 13628
rect 18256 13572 18312 13628
rect 18312 13572 18316 13628
rect 18252 13568 18316 13572
rect 18332 13628 18396 13632
rect 18332 13572 18336 13628
rect 18336 13572 18392 13628
rect 18392 13572 18396 13628
rect 18332 13568 18396 13572
rect 18412 13628 18476 13632
rect 18412 13572 18416 13628
rect 18416 13572 18472 13628
rect 18472 13572 18476 13628
rect 18412 13568 18476 13572
rect 18492 13628 18556 13632
rect 18492 13572 18496 13628
rect 18496 13572 18552 13628
rect 18552 13572 18556 13628
rect 18492 13568 18556 13572
rect 21252 13628 21316 13632
rect 21252 13572 21256 13628
rect 21256 13572 21312 13628
rect 21312 13572 21316 13628
rect 21252 13568 21316 13572
rect 21332 13628 21396 13632
rect 21332 13572 21336 13628
rect 21336 13572 21392 13628
rect 21392 13572 21396 13628
rect 21332 13568 21396 13572
rect 21412 13628 21476 13632
rect 21412 13572 21416 13628
rect 21416 13572 21472 13628
rect 21472 13572 21476 13628
rect 21412 13568 21476 13572
rect 21492 13628 21556 13632
rect 21492 13572 21496 13628
rect 21496 13572 21552 13628
rect 21552 13572 21556 13628
rect 21492 13568 21556 13572
rect 24252 13628 24316 13632
rect 24252 13572 24256 13628
rect 24256 13572 24312 13628
rect 24312 13572 24316 13628
rect 24252 13568 24316 13572
rect 24332 13628 24396 13632
rect 24332 13572 24336 13628
rect 24336 13572 24392 13628
rect 24392 13572 24396 13628
rect 24332 13568 24396 13572
rect 24412 13628 24476 13632
rect 24412 13572 24416 13628
rect 24416 13572 24472 13628
rect 24472 13572 24476 13628
rect 24412 13568 24476 13572
rect 24492 13628 24556 13632
rect 24492 13572 24496 13628
rect 24496 13572 24552 13628
rect 24552 13572 24556 13628
rect 24492 13568 24556 13572
rect 27252 13628 27316 13632
rect 27252 13572 27256 13628
rect 27256 13572 27312 13628
rect 27312 13572 27316 13628
rect 27252 13568 27316 13572
rect 27332 13628 27396 13632
rect 27332 13572 27336 13628
rect 27336 13572 27392 13628
rect 27392 13572 27396 13628
rect 27332 13568 27396 13572
rect 27412 13628 27476 13632
rect 27412 13572 27416 13628
rect 27416 13572 27472 13628
rect 27472 13572 27476 13628
rect 27412 13568 27476 13572
rect 27492 13628 27556 13632
rect 27492 13572 27496 13628
rect 27496 13572 27552 13628
rect 27552 13572 27556 13628
rect 27492 13568 27556 13572
rect 1752 13084 1816 13088
rect 1752 13028 1756 13084
rect 1756 13028 1812 13084
rect 1812 13028 1816 13084
rect 1752 13024 1816 13028
rect 1832 13084 1896 13088
rect 1832 13028 1836 13084
rect 1836 13028 1892 13084
rect 1892 13028 1896 13084
rect 1832 13024 1896 13028
rect 1912 13084 1976 13088
rect 1912 13028 1916 13084
rect 1916 13028 1972 13084
rect 1972 13028 1976 13084
rect 1912 13024 1976 13028
rect 1992 13084 2056 13088
rect 1992 13028 1996 13084
rect 1996 13028 2052 13084
rect 2052 13028 2056 13084
rect 1992 13024 2056 13028
rect 4752 13084 4816 13088
rect 4752 13028 4756 13084
rect 4756 13028 4812 13084
rect 4812 13028 4816 13084
rect 4752 13024 4816 13028
rect 4832 13084 4896 13088
rect 4832 13028 4836 13084
rect 4836 13028 4892 13084
rect 4892 13028 4896 13084
rect 4832 13024 4896 13028
rect 4912 13084 4976 13088
rect 4912 13028 4916 13084
rect 4916 13028 4972 13084
rect 4972 13028 4976 13084
rect 4912 13024 4976 13028
rect 4992 13084 5056 13088
rect 4992 13028 4996 13084
rect 4996 13028 5052 13084
rect 5052 13028 5056 13084
rect 4992 13024 5056 13028
rect 7752 13084 7816 13088
rect 7752 13028 7756 13084
rect 7756 13028 7812 13084
rect 7812 13028 7816 13084
rect 7752 13024 7816 13028
rect 7832 13084 7896 13088
rect 7832 13028 7836 13084
rect 7836 13028 7892 13084
rect 7892 13028 7896 13084
rect 7832 13024 7896 13028
rect 7912 13084 7976 13088
rect 7912 13028 7916 13084
rect 7916 13028 7972 13084
rect 7972 13028 7976 13084
rect 7912 13024 7976 13028
rect 7992 13084 8056 13088
rect 7992 13028 7996 13084
rect 7996 13028 8052 13084
rect 8052 13028 8056 13084
rect 7992 13024 8056 13028
rect 10752 13084 10816 13088
rect 10752 13028 10756 13084
rect 10756 13028 10812 13084
rect 10812 13028 10816 13084
rect 10752 13024 10816 13028
rect 10832 13084 10896 13088
rect 10832 13028 10836 13084
rect 10836 13028 10892 13084
rect 10892 13028 10896 13084
rect 10832 13024 10896 13028
rect 10912 13084 10976 13088
rect 10912 13028 10916 13084
rect 10916 13028 10972 13084
rect 10972 13028 10976 13084
rect 10912 13024 10976 13028
rect 10992 13084 11056 13088
rect 10992 13028 10996 13084
rect 10996 13028 11052 13084
rect 11052 13028 11056 13084
rect 10992 13024 11056 13028
rect 13752 13084 13816 13088
rect 13752 13028 13756 13084
rect 13756 13028 13812 13084
rect 13812 13028 13816 13084
rect 13752 13024 13816 13028
rect 13832 13084 13896 13088
rect 13832 13028 13836 13084
rect 13836 13028 13892 13084
rect 13892 13028 13896 13084
rect 13832 13024 13896 13028
rect 13912 13084 13976 13088
rect 13912 13028 13916 13084
rect 13916 13028 13972 13084
rect 13972 13028 13976 13084
rect 13912 13024 13976 13028
rect 13992 13084 14056 13088
rect 13992 13028 13996 13084
rect 13996 13028 14052 13084
rect 14052 13028 14056 13084
rect 13992 13024 14056 13028
rect 16752 13084 16816 13088
rect 16752 13028 16756 13084
rect 16756 13028 16812 13084
rect 16812 13028 16816 13084
rect 16752 13024 16816 13028
rect 16832 13084 16896 13088
rect 16832 13028 16836 13084
rect 16836 13028 16892 13084
rect 16892 13028 16896 13084
rect 16832 13024 16896 13028
rect 16912 13084 16976 13088
rect 16912 13028 16916 13084
rect 16916 13028 16972 13084
rect 16972 13028 16976 13084
rect 16912 13024 16976 13028
rect 16992 13084 17056 13088
rect 16992 13028 16996 13084
rect 16996 13028 17052 13084
rect 17052 13028 17056 13084
rect 16992 13024 17056 13028
rect 19752 13084 19816 13088
rect 19752 13028 19756 13084
rect 19756 13028 19812 13084
rect 19812 13028 19816 13084
rect 19752 13024 19816 13028
rect 19832 13084 19896 13088
rect 19832 13028 19836 13084
rect 19836 13028 19892 13084
rect 19892 13028 19896 13084
rect 19832 13024 19896 13028
rect 19912 13084 19976 13088
rect 19912 13028 19916 13084
rect 19916 13028 19972 13084
rect 19972 13028 19976 13084
rect 19912 13024 19976 13028
rect 19992 13084 20056 13088
rect 19992 13028 19996 13084
rect 19996 13028 20052 13084
rect 20052 13028 20056 13084
rect 19992 13024 20056 13028
rect 22752 13084 22816 13088
rect 22752 13028 22756 13084
rect 22756 13028 22812 13084
rect 22812 13028 22816 13084
rect 22752 13024 22816 13028
rect 22832 13084 22896 13088
rect 22832 13028 22836 13084
rect 22836 13028 22892 13084
rect 22892 13028 22896 13084
rect 22832 13024 22896 13028
rect 22912 13084 22976 13088
rect 22912 13028 22916 13084
rect 22916 13028 22972 13084
rect 22972 13028 22976 13084
rect 22912 13024 22976 13028
rect 22992 13084 23056 13088
rect 22992 13028 22996 13084
rect 22996 13028 23052 13084
rect 23052 13028 23056 13084
rect 22992 13024 23056 13028
rect 25752 13084 25816 13088
rect 25752 13028 25756 13084
rect 25756 13028 25812 13084
rect 25812 13028 25816 13084
rect 25752 13024 25816 13028
rect 25832 13084 25896 13088
rect 25832 13028 25836 13084
rect 25836 13028 25892 13084
rect 25892 13028 25896 13084
rect 25832 13024 25896 13028
rect 25912 13084 25976 13088
rect 25912 13028 25916 13084
rect 25916 13028 25972 13084
rect 25972 13028 25976 13084
rect 25912 13024 25976 13028
rect 25992 13084 26056 13088
rect 25992 13028 25996 13084
rect 25996 13028 26052 13084
rect 26052 13028 26056 13084
rect 25992 13024 26056 13028
rect 3252 12540 3316 12544
rect 3252 12484 3256 12540
rect 3256 12484 3312 12540
rect 3312 12484 3316 12540
rect 3252 12480 3316 12484
rect 3332 12540 3396 12544
rect 3332 12484 3336 12540
rect 3336 12484 3392 12540
rect 3392 12484 3396 12540
rect 3332 12480 3396 12484
rect 3412 12540 3476 12544
rect 3412 12484 3416 12540
rect 3416 12484 3472 12540
rect 3472 12484 3476 12540
rect 3412 12480 3476 12484
rect 3492 12540 3556 12544
rect 3492 12484 3496 12540
rect 3496 12484 3552 12540
rect 3552 12484 3556 12540
rect 3492 12480 3556 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 6412 12540 6476 12544
rect 6412 12484 6416 12540
rect 6416 12484 6472 12540
rect 6472 12484 6476 12540
rect 6412 12480 6476 12484
rect 6492 12540 6556 12544
rect 6492 12484 6496 12540
rect 6496 12484 6552 12540
rect 6552 12484 6556 12540
rect 6492 12480 6556 12484
rect 9252 12540 9316 12544
rect 9252 12484 9256 12540
rect 9256 12484 9312 12540
rect 9312 12484 9316 12540
rect 9252 12480 9316 12484
rect 9332 12540 9396 12544
rect 9332 12484 9336 12540
rect 9336 12484 9392 12540
rect 9392 12484 9396 12540
rect 9332 12480 9396 12484
rect 9412 12540 9476 12544
rect 9412 12484 9416 12540
rect 9416 12484 9472 12540
rect 9472 12484 9476 12540
rect 9412 12480 9476 12484
rect 9492 12540 9556 12544
rect 9492 12484 9496 12540
rect 9496 12484 9552 12540
rect 9552 12484 9556 12540
rect 9492 12480 9556 12484
rect 12252 12540 12316 12544
rect 12252 12484 12256 12540
rect 12256 12484 12312 12540
rect 12312 12484 12316 12540
rect 12252 12480 12316 12484
rect 12332 12540 12396 12544
rect 12332 12484 12336 12540
rect 12336 12484 12392 12540
rect 12392 12484 12396 12540
rect 12332 12480 12396 12484
rect 12412 12540 12476 12544
rect 12412 12484 12416 12540
rect 12416 12484 12472 12540
rect 12472 12484 12476 12540
rect 12412 12480 12476 12484
rect 12492 12540 12556 12544
rect 12492 12484 12496 12540
rect 12496 12484 12552 12540
rect 12552 12484 12556 12540
rect 12492 12480 12556 12484
rect 15252 12540 15316 12544
rect 15252 12484 15256 12540
rect 15256 12484 15312 12540
rect 15312 12484 15316 12540
rect 15252 12480 15316 12484
rect 15332 12540 15396 12544
rect 15332 12484 15336 12540
rect 15336 12484 15392 12540
rect 15392 12484 15396 12540
rect 15332 12480 15396 12484
rect 15412 12540 15476 12544
rect 15412 12484 15416 12540
rect 15416 12484 15472 12540
rect 15472 12484 15476 12540
rect 15412 12480 15476 12484
rect 15492 12540 15556 12544
rect 15492 12484 15496 12540
rect 15496 12484 15552 12540
rect 15552 12484 15556 12540
rect 15492 12480 15556 12484
rect 18252 12540 18316 12544
rect 18252 12484 18256 12540
rect 18256 12484 18312 12540
rect 18312 12484 18316 12540
rect 18252 12480 18316 12484
rect 18332 12540 18396 12544
rect 18332 12484 18336 12540
rect 18336 12484 18392 12540
rect 18392 12484 18396 12540
rect 18332 12480 18396 12484
rect 18412 12540 18476 12544
rect 18412 12484 18416 12540
rect 18416 12484 18472 12540
rect 18472 12484 18476 12540
rect 18412 12480 18476 12484
rect 18492 12540 18556 12544
rect 18492 12484 18496 12540
rect 18496 12484 18552 12540
rect 18552 12484 18556 12540
rect 18492 12480 18556 12484
rect 21252 12540 21316 12544
rect 21252 12484 21256 12540
rect 21256 12484 21312 12540
rect 21312 12484 21316 12540
rect 21252 12480 21316 12484
rect 21332 12540 21396 12544
rect 21332 12484 21336 12540
rect 21336 12484 21392 12540
rect 21392 12484 21396 12540
rect 21332 12480 21396 12484
rect 21412 12540 21476 12544
rect 21412 12484 21416 12540
rect 21416 12484 21472 12540
rect 21472 12484 21476 12540
rect 21412 12480 21476 12484
rect 21492 12540 21556 12544
rect 21492 12484 21496 12540
rect 21496 12484 21552 12540
rect 21552 12484 21556 12540
rect 21492 12480 21556 12484
rect 24252 12540 24316 12544
rect 24252 12484 24256 12540
rect 24256 12484 24312 12540
rect 24312 12484 24316 12540
rect 24252 12480 24316 12484
rect 24332 12540 24396 12544
rect 24332 12484 24336 12540
rect 24336 12484 24392 12540
rect 24392 12484 24396 12540
rect 24332 12480 24396 12484
rect 24412 12540 24476 12544
rect 24412 12484 24416 12540
rect 24416 12484 24472 12540
rect 24472 12484 24476 12540
rect 24412 12480 24476 12484
rect 24492 12540 24556 12544
rect 24492 12484 24496 12540
rect 24496 12484 24552 12540
rect 24552 12484 24556 12540
rect 24492 12480 24556 12484
rect 27252 12540 27316 12544
rect 27252 12484 27256 12540
rect 27256 12484 27312 12540
rect 27312 12484 27316 12540
rect 27252 12480 27316 12484
rect 27332 12540 27396 12544
rect 27332 12484 27336 12540
rect 27336 12484 27392 12540
rect 27392 12484 27396 12540
rect 27332 12480 27396 12484
rect 27412 12540 27476 12544
rect 27412 12484 27416 12540
rect 27416 12484 27472 12540
rect 27472 12484 27476 12540
rect 27412 12480 27476 12484
rect 27492 12540 27556 12544
rect 27492 12484 27496 12540
rect 27496 12484 27552 12540
rect 27552 12484 27556 12540
rect 27492 12480 27556 12484
rect 1752 11996 1816 12000
rect 1752 11940 1756 11996
rect 1756 11940 1812 11996
rect 1812 11940 1816 11996
rect 1752 11936 1816 11940
rect 1832 11996 1896 12000
rect 1832 11940 1836 11996
rect 1836 11940 1892 11996
rect 1892 11940 1896 11996
rect 1832 11936 1896 11940
rect 1912 11996 1976 12000
rect 1912 11940 1916 11996
rect 1916 11940 1972 11996
rect 1972 11940 1976 11996
rect 1912 11936 1976 11940
rect 1992 11996 2056 12000
rect 1992 11940 1996 11996
rect 1996 11940 2052 11996
rect 2052 11940 2056 11996
rect 1992 11936 2056 11940
rect 4752 11996 4816 12000
rect 4752 11940 4756 11996
rect 4756 11940 4812 11996
rect 4812 11940 4816 11996
rect 4752 11936 4816 11940
rect 4832 11996 4896 12000
rect 4832 11940 4836 11996
rect 4836 11940 4892 11996
rect 4892 11940 4896 11996
rect 4832 11936 4896 11940
rect 4912 11996 4976 12000
rect 4912 11940 4916 11996
rect 4916 11940 4972 11996
rect 4972 11940 4976 11996
rect 4912 11936 4976 11940
rect 4992 11996 5056 12000
rect 4992 11940 4996 11996
rect 4996 11940 5052 11996
rect 5052 11940 5056 11996
rect 4992 11936 5056 11940
rect 7752 11996 7816 12000
rect 7752 11940 7756 11996
rect 7756 11940 7812 11996
rect 7812 11940 7816 11996
rect 7752 11936 7816 11940
rect 7832 11996 7896 12000
rect 7832 11940 7836 11996
rect 7836 11940 7892 11996
rect 7892 11940 7896 11996
rect 7832 11936 7896 11940
rect 7912 11996 7976 12000
rect 7912 11940 7916 11996
rect 7916 11940 7972 11996
rect 7972 11940 7976 11996
rect 7912 11936 7976 11940
rect 7992 11996 8056 12000
rect 7992 11940 7996 11996
rect 7996 11940 8052 11996
rect 8052 11940 8056 11996
rect 7992 11936 8056 11940
rect 10752 11996 10816 12000
rect 10752 11940 10756 11996
rect 10756 11940 10812 11996
rect 10812 11940 10816 11996
rect 10752 11936 10816 11940
rect 10832 11996 10896 12000
rect 10832 11940 10836 11996
rect 10836 11940 10892 11996
rect 10892 11940 10896 11996
rect 10832 11936 10896 11940
rect 10912 11996 10976 12000
rect 10912 11940 10916 11996
rect 10916 11940 10972 11996
rect 10972 11940 10976 11996
rect 10912 11936 10976 11940
rect 10992 11996 11056 12000
rect 10992 11940 10996 11996
rect 10996 11940 11052 11996
rect 11052 11940 11056 11996
rect 10992 11936 11056 11940
rect 13752 11996 13816 12000
rect 13752 11940 13756 11996
rect 13756 11940 13812 11996
rect 13812 11940 13816 11996
rect 13752 11936 13816 11940
rect 13832 11996 13896 12000
rect 13832 11940 13836 11996
rect 13836 11940 13892 11996
rect 13892 11940 13896 11996
rect 13832 11936 13896 11940
rect 13912 11996 13976 12000
rect 13912 11940 13916 11996
rect 13916 11940 13972 11996
rect 13972 11940 13976 11996
rect 13912 11936 13976 11940
rect 13992 11996 14056 12000
rect 13992 11940 13996 11996
rect 13996 11940 14052 11996
rect 14052 11940 14056 11996
rect 13992 11936 14056 11940
rect 16752 11996 16816 12000
rect 16752 11940 16756 11996
rect 16756 11940 16812 11996
rect 16812 11940 16816 11996
rect 16752 11936 16816 11940
rect 16832 11996 16896 12000
rect 16832 11940 16836 11996
rect 16836 11940 16892 11996
rect 16892 11940 16896 11996
rect 16832 11936 16896 11940
rect 16912 11996 16976 12000
rect 16912 11940 16916 11996
rect 16916 11940 16972 11996
rect 16972 11940 16976 11996
rect 16912 11936 16976 11940
rect 16992 11996 17056 12000
rect 16992 11940 16996 11996
rect 16996 11940 17052 11996
rect 17052 11940 17056 11996
rect 16992 11936 17056 11940
rect 19752 11996 19816 12000
rect 19752 11940 19756 11996
rect 19756 11940 19812 11996
rect 19812 11940 19816 11996
rect 19752 11936 19816 11940
rect 19832 11996 19896 12000
rect 19832 11940 19836 11996
rect 19836 11940 19892 11996
rect 19892 11940 19896 11996
rect 19832 11936 19896 11940
rect 19912 11996 19976 12000
rect 19912 11940 19916 11996
rect 19916 11940 19972 11996
rect 19972 11940 19976 11996
rect 19912 11936 19976 11940
rect 19992 11996 20056 12000
rect 19992 11940 19996 11996
rect 19996 11940 20052 11996
rect 20052 11940 20056 11996
rect 19992 11936 20056 11940
rect 22752 11996 22816 12000
rect 22752 11940 22756 11996
rect 22756 11940 22812 11996
rect 22812 11940 22816 11996
rect 22752 11936 22816 11940
rect 22832 11996 22896 12000
rect 22832 11940 22836 11996
rect 22836 11940 22892 11996
rect 22892 11940 22896 11996
rect 22832 11936 22896 11940
rect 22912 11996 22976 12000
rect 22912 11940 22916 11996
rect 22916 11940 22972 11996
rect 22972 11940 22976 11996
rect 22912 11936 22976 11940
rect 22992 11996 23056 12000
rect 22992 11940 22996 11996
rect 22996 11940 23052 11996
rect 23052 11940 23056 11996
rect 22992 11936 23056 11940
rect 25752 11996 25816 12000
rect 25752 11940 25756 11996
rect 25756 11940 25812 11996
rect 25812 11940 25816 11996
rect 25752 11936 25816 11940
rect 25832 11996 25896 12000
rect 25832 11940 25836 11996
rect 25836 11940 25892 11996
rect 25892 11940 25896 11996
rect 25832 11936 25896 11940
rect 25912 11996 25976 12000
rect 25912 11940 25916 11996
rect 25916 11940 25972 11996
rect 25972 11940 25976 11996
rect 25912 11936 25976 11940
rect 25992 11996 26056 12000
rect 25992 11940 25996 11996
rect 25996 11940 26052 11996
rect 26052 11940 26056 11996
rect 25992 11936 26056 11940
rect 3252 11452 3316 11456
rect 3252 11396 3256 11452
rect 3256 11396 3312 11452
rect 3312 11396 3316 11452
rect 3252 11392 3316 11396
rect 3332 11452 3396 11456
rect 3332 11396 3336 11452
rect 3336 11396 3392 11452
rect 3392 11396 3396 11452
rect 3332 11392 3396 11396
rect 3412 11452 3476 11456
rect 3412 11396 3416 11452
rect 3416 11396 3472 11452
rect 3472 11396 3476 11452
rect 3412 11392 3476 11396
rect 3492 11452 3556 11456
rect 3492 11396 3496 11452
rect 3496 11396 3552 11452
rect 3552 11396 3556 11452
rect 3492 11392 3556 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 6412 11452 6476 11456
rect 6412 11396 6416 11452
rect 6416 11396 6472 11452
rect 6472 11396 6476 11452
rect 6412 11392 6476 11396
rect 6492 11452 6556 11456
rect 6492 11396 6496 11452
rect 6496 11396 6552 11452
rect 6552 11396 6556 11452
rect 6492 11392 6556 11396
rect 9252 11452 9316 11456
rect 9252 11396 9256 11452
rect 9256 11396 9312 11452
rect 9312 11396 9316 11452
rect 9252 11392 9316 11396
rect 9332 11452 9396 11456
rect 9332 11396 9336 11452
rect 9336 11396 9392 11452
rect 9392 11396 9396 11452
rect 9332 11392 9396 11396
rect 9412 11452 9476 11456
rect 9412 11396 9416 11452
rect 9416 11396 9472 11452
rect 9472 11396 9476 11452
rect 9412 11392 9476 11396
rect 9492 11452 9556 11456
rect 9492 11396 9496 11452
rect 9496 11396 9552 11452
rect 9552 11396 9556 11452
rect 9492 11392 9556 11396
rect 12252 11452 12316 11456
rect 12252 11396 12256 11452
rect 12256 11396 12312 11452
rect 12312 11396 12316 11452
rect 12252 11392 12316 11396
rect 12332 11452 12396 11456
rect 12332 11396 12336 11452
rect 12336 11396 12392 11452
rect 12392 11396 12396 11452
rect 12332 11392 12396 11396
rect 12412 11452 12476 11456
rect 12412 11396 12416 11452
rect 12416 11396 12472 11452
rect 12472 11396 12476 11452
rect 12412 11392 12476 11396
rect 12492 11452 12556 11456
rect 12492 11396 12496 11452
rect 12496 11396 12552 11452
rect 12552 11396 12556 11452
rect 12492 11392 12556 11396
rect 15252 11452 15316 11456
rect 15252 11396 15256 11452
rect 15256 11396 15312 11452
rect 15312 11396 15316 11452
rect 15252 11392 15316 11396
rect 15332 11452 15396 11456
rect 15332 11396 15336 11452
rect 15336 11396 15392 11452
rect 15392 11396 15396 11452
rect 15332 11392 15396 11396
rect 15412 11452 15476 11456
rect 15412 11396 15416 11452
rect 15416 11396 15472 11452
rect 15472 11396 15476 11452
rect 15412 11392 15476 11396
rect 15492 11452 15556 11456
rect 15492 11396 15496 11452
rect 15496 11396 15552 11452
rect 15552 11396 15556 11452
rect 15492 11392 15556 11396
rect 18252 11452 18316 11456
rect 18252 11396 18256 11452
rect 18256 11396 18312 11452
rect 18312 11396 18316 11452
rect 18252 11392 18316 11396
rect 18332 11452 18396 11456
rect 18332 11396 18336 11452
rect 18336 11396 18392 11452
rect 18392 11396 18396 11452
rect 18332 11392 18396 11396
rect 18412 11452 18476 11456
rect 18412 11396 18416 11452
rect 18416 11396 18472 11452
rect 18472 11396 18476 11452
rect 18412 11392 18476 11396
rect 18492 11452 18556 11456
rect 18492 11396 18496 11452
rect 18496 11396 18552 11452
rect 18552 11396 18556 11452
rect 18492 11392 18556 11396
rect 21252 11452 21316 11456
rect 21252 11396 21256 11452
rect 21256 11396 21312 11452
rect 21312 11396 21316 11452
rect 21252 11392 21316 11396
rect 21332 11452 21396 11456
rect 21332 11396 21336 11452
rect 21336 11396 21392 11452
rect 21392 11396 21396 11452
rect 21332 11392 21396 11396
rect 21412 11452 21476 11456
rect 21412 11396 21416 11452
rect 21416 11396 21472 11452
rect 21472 11396 21476 11452
rect 21412 11392 21476 11396
rect 21492 11452 21556 11456
rect 21492 11396 21496 11452
rect 21496 11396 21552 11452
rect 21552 11396 21556 11452
rect 21492 11392 21556 11396
rect 24252 11452 24316 11456
rect 24252 11396 24256 11452
rect 24256 11396 24312 11452
rect 24312 11396 24316 11452
rect 24252 11392 24316 11396
rect 24332 11452 24396 11456
rect 24332 11396 24336 11452
rect 24336 11396 24392 11452
rect 24392 11396 24396 11452
rect 24332 11392 24396 11396
rect 24412 11452 24476 11456
rect 24412 11396 24416 11452
rect 24416 11396 24472 11452
rect 24472 11396 24476 11452
rect 24412 11392 24476 11396
rect 24492 11452 24556 11456
rect 24492 11396 24496 11452
rect 24496 11396 24552 11452
rect 24552 11396 24556 11452
rect 24492 11392 24556 11396
rect 27252 11452 27316 11456
rect 27252 11396 27256 11452
rect 27256 11396 27312 11452
rect 27312 11396 27316 11452
rect 27252 11392 27316 11396
rect 27332 11452 27396 11456
rect 27332 11396 27336 11452
rect 27336 11396 27392 11452
rect 27392 11396 27396 11452
rect 27332 11392 27396 11396
rect 27412 11452 27476 11456
rect 27412 11396 27416 11452
rect 27416 11396 27472 11452
rect 27472 11396 27476 11452
rect 27412 11392 27476 11396
rect 27492 11452 27556 11456
rect 27492 11396 27496 11452
rect 27496 11396 27552 11452
rect 27552 11396 27556 11452
rect 27492 11392 27556 11396
rect 1752 10908 1816 10912
rect 1752 10852 1756 10908
rect 1756 10852 1812 10908
rect 1812 10852 1816 10908
rect 1752 10848 1816 10852
rect 1832 10908 1896 10912
rect 1832 10852 1836 10908
rect 1836 10852 1892 10908
rect 1892 10852 1896 10908
rect 1832 10848 1896 10852
rect 1912 10908 1976 10912
rect 1912 10852 1916 10908
rect 1916 10852 1972 10908
rect 1972 10852 1976 10908
rect 1912 10848 1976 10852
rect 1992 10908 2056 10912
rect 1992 10852 1996 10908
rect 1996 10852 2052 10908
rect 2052 10852 2056 10908
rect 1992 10848 2056 10852
rect 4752 10908 4816 10912
rect 4752 10852 4756 10908
rect 4756 10852 4812 10908
rect 4812 10852 4816 10908
rect 4752 10848 4816 10852
rect 4832 10908 4896 10912
rect 4832 10852 4836 10908
rect 4836 10852 4892 10908
rect 4892 10852 4896 10908
rect 4832 10848 4896 10852
rect 4912 10908 4976 10912
rect 4912 10852 4916 10908
rect 4916 10852 4972 10908
rect 4972 10852 4976 10908
rect 4912 10848 4976 10852
rect 4992 10908 5056 10912
rect 4992 10852 4996 10908
rect 4996 10852 5052 10908
rect 5052 10852 5056 10908
rect 4992 10848 5056 10852
rect 7752 10908 7816 10912
rect 7752 10852 7756 10908
rect 7756 10852 7812 10908
rect 7812 10852 7816 10908
rect 7752 10848 7816 10852
rect 7832 10908 7896 10912
rect 7832 10852 7836 10908
rect 7836 10852 7892 10908
rect 7892 10852 7896 10908
rect 7832 10848 7896 10852
rect 7912 10908 7976 10912
rect 7912 10852 7916 10908
rect 7916 10852 7972 10908
rect 7972 10852 7976 10908
rect 7912 10848 7976 10852
rect 7992 10908 8056 10912
rect 7992 10852 7996 10908
rect 7996 10852 8052 10908
rect 8052 10852 8056 10908
rect 7992 10848 8056 10852
rect 10752 10908 10816 10912
rect 10752 10852 10756 10908
rect 10756 10852 10812 10908
rect 10812 10852 10816 10908
rect 10752 10848 10816 10852
rect 10832 10908 10896 10912
rect 10832 10852 10836 10908
rect 10836 10852 10892 10908
rect 10892 10852 10896 10908
rect 10832 10848 10896 10852
rect 10912 10908 10976 10912
rect 10912 10852 10916 10908
rect 10916 10852 10972 10908
rect 10972 10852 10976 10908
rect 10912 10848 10976 10852
rect 10992 10908 11056 10912
rect 10992 10852 10996 10908
rect 10996 10852 11052 10908
rect 11052 10852 11056 10908
rect 10992 10848 11056 10852
rect 13752 10908 13816 10912
rect 13752 10852 13756 10908
rect 13756 10852 13812 10908
rect 13812 10852 13816 10908
rect 13752 10848 13816 10852
rect 13832 10908 13896 10912
rect 13832 10852 13836 10908
rect 13836 10852 13892 10908
rect 13892 10852 13896 10908
rect 13832 10848 13896 10852
rect 13912 10908 13976 10912
rect 13912 10852 13916 10908
rect 13916 10852 13972 10908
rect 13972 10852 13976 10908
rect 13912 10848 13976 10852
rect 13992 10908 14056 10912
rect 13992 10852 13996 10908
rect 13996 10852 14052 10908
rect 14052 10852 14056 10908
rect 13992 10848 14056 10852
rect 16752 10908 16816 10912
rect 16752 10852 16756 10908
rect 16756 10852 16812 10908
rect 16812 10852 16816 10908
rect 16752 10848 16816 10852
rect 16832 10908 16896 10912
rect 16832 10852 16836 10908
rect 16836 10852 16892 10908
rect 16892 10852 16896 10908
rect 16832 10848 16896 10852
rect 16912 10908 16976 10912
rect 16912 10852 16916 10908
rect 16916 10852 16972 10908
rect 16972 10852 16976 10908
rect 16912 10848 16976 10852
rect 16992 10908 17056 10912
rect 16992 10852 16996 10908
rect 16996 10852 17052 10908
rect 17052 10852 17056 10908
rect 16992 10848 17056 10852
rect 19752 10908 19816 10912
rect 19752 10852 19756 10908
rect 19756 10852 19812 10908
rect 19812 10852 19816 10908
rect 19752 10848 19816 10852
rect 19832 10908 19896 10912
rect 19832 10852 19836 10908
rect 19836 10852 19892 10908
rect 19892 10852 19896 10908
rect 19832 10848 19896 10852
rect 19912 10908 19976 10912
rect 19912 10852 19916 10908
rect 19916 10852 19972 10908
rect 19972 10852 19976 10908
rect 19912 10848 19976 10852
rect 19992 10908 20056 10912
rect 19992 10852 19996 10908
rect 19996 10852 20052 10908
rect 20052 10852 20056 10908
rect 19992 10848 20056 10852
rect 22752 10908 22816 10912
rect 22752 10852 22756 10908
rect 22756 10852 22812 10908
rect 22812 10852 22816 10908
rect 22752 10848 22816 10852
rect 22832 10908 22896 10912
rect 22832 10852 22836 10908
rect 22836 10852 22892 10908
rect 22892 10852 22896 10908
rect 22832 10848 22896 10852
rect 22912 10908 22976 10912
rect 22912 10852 22916 10908
rect 22916 10852 22972 10908
rect 22972 10852 22976 10908
rect 22912 10848 22976 10852
rect 22992 10908 23056 10912
rect 22992 10852 22996 10908
rect 22996 10852 23052 10908
rect 23052 10852 23056 10908
rect 22992 10848 23056 10852
rect 25752 10908 25816 10912
rect 25752 10852 25756 10908
rect 25756 10852 25812 10908
rect 25812 10852 25816 10908
rect 25752 10848 25816 10852
rect 25832 10908 25896 10912
rect 25832 10852 25836 10908
rect 25836 10852 25892 10908
rect 25892 10852 25896 10908
rect 25832 10848 25896 10852
rect 25912 10908 25976 10912
rect 25912 10852 25916 10908
rect 25916 10852 25972 10908
rect 25972 10852 25976 10908
rect 25912 10848 25976 10852
rect 25992 10908 26056 10912
rect 25992 10852 25996 10908
rect 25996 10852 26052 10908
rect 26052 10852 26056 10908
rect 25992 10848 26056 10852
rect 3252 10364 3316 10368
rect 3252 10308 3256 10364
rect 3256 10308 3312 10364
rect 3312 10308 3316 10364
rect 3252 10304 3316 10308
rect 3332 10364 3396 10368
rect 3332 10308 3336 10364
rect 3336 10308 3392 10364
rect 3392 10308 3396 10364
rect 3332 10304 3396 10308
rect 3412 10364 3476 10368
rect 3412 10308 3416 10364
rect 3416 10308 3472 10364
rect 3472 10308 3476 10364
rect 3412 10304 3476 10308
rect 3492 10364 3556 10368
rect 3492 10308 3496 10364
rect 3496 10308 3552 10364
rect 3552 10308 3556 10364
rect 3492 10304 3556 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 6412 10364 6476 10368
rect 6412 10308 6416 10364
rect 6416 10308 6472 10364
rect 6472 10308 6476 10364
rect 6412 10304 6476 10308
rect 6492 10364 6556 10368
rect 6492 10308 6496 10364
rect 6496 10308 6552 10364
rect 6552 10308 6556 10364
rect 6492 10304 6556 10308
rect 9252 10364 9316 10368
rect 9252 10308 9256 10364
rect 9256 10308 9312 10364
rect 9312 10308 9316 10364
rect 9252 10304 9316 10308
rect 9332 10364 9396 10368
rect 9332 10308 9336 10364
rect 9336 10308 9392 10364
rect 9392 10308 9396 10364
rect 9332 10304 9396 10308
rect 9412 10364 9476 10368
rect 9412 10308 9416 10364
rect 9416 10308 9472 10364
rect 9472 10308 9476 10364
rect 9412 10304 9476 10308
rect 9492 10364 9556 10368
rect 9492 10308 9496 10364
rect 9496 10308 9552 10364
rect 9552 10308 9556 10364
rect 9492 10304 9556 10308
rect 12252 10364 12316 10368
rect 12252 10308 12256 10364
rect 12256 10308 12312 10364
rect 12312 10308 12316 10364
rect 12252 10304 12316 10308
rect 12332 10364 12396 10368
rect 12332 10308 12336 10364
rect 12336 10308 12392 10364
rect 12392 10308 12396 10364
rect 12332 10304 12396 10308
rect 12412 10364 12476 10368
rect 12412 10308 12416 10364
rect 12416 10308 12472 10364
rect 12472 10308 12476 10364
rect 12412 10304 12476 10308
rect 12492 10364 12556 10368
rect 12492 10308 12496 10364
rect 12496 10308 12552 10364
rect 12552 10308 12556 10364
rect 12492 10304 12556 10308
rect 15252 10364 15316 10368
rect 15252 10308 15256 10364
rect 15256 10308 15312 10364
rect 15312 10308 15316 10364
rect 15252 10304 15316 10308
rect 15332 10364 15396 10368
rect 15332 10308 15336 10364
rect 15336 10308 15392 10364
rect 15392 10308 15396 10364
rect 15332 10304 15396 10308
rect 15412 10364 15476 10368
rect 15412 10308 15416 10364
rect 15416 10308 15472 10364
rect 15472 10308 15476 10364
rect 15412 10304 15476 10308
rect 15492 10364 15556 10368
rect 15492 10308 15496 10364
rect 15496 10308 15552 10364
rect 15552 10308 15556 10364
rect 15492 10304 15556 10308
rect 18252 10364 18316 10368
rect 18252 10308 18256 10364
rect 18256 10308 18312 10364
rect 18312 10308 18316 10364
rect 18252 10304 18316 10308
rect 18332 10364 18396 10368
rect 18332 10308 18336 10364
rect 18336 10308 18392 10364
rect 18392 10308 18396 10364
rect 18332 10304 18396 10308
rect 18412 10364 18476 10368
rect 18412 10308 18416 10364
rect 18416 10308 18472 10364
rect 18472 10308 18476 10364
rect 18412 10304 18476 10308
rect 18492 10364 18556 10368
rect 18492 10308 18496 10364
rect 18496 10308 18552 10364
rect 18552 10308 18556 10364
rect 18492 10304 18556 10308
rect 21252 10364 21316 10368
rect 21252 10308 21256 10364
rect 21256 10308 21312 10364
rect 21312 10308 21316 10364
rect 21252 10304 21316 10308
rect 21332 10364 21396 10368
rect 21332 10308 21336 10364
rect 21336 10308 21392 10364
rect 21392 10308 21396 10364
rect 21332 10304 21396 10308
rect 21412 10364 21476 10368
rect 21412 10308 21416 10364
rect 21416 10308 21472 10364
rect 21472 10308 21476 10364
rect 21412 10304 21476 10308
rect 21492 10364 21556 10368
rect 21492 10308 21496 10364
rect 21496 10308 21552 10364
rect 21552 10308 21556 10364
rect 21492 10304 21556 10308
rect 24252 10364 24316 10368
rect 24252 10308 24256 10364
rect 24256 10308 24312 10364
rect 24312 10308 24316 10364
rect 24252 10304 24316 10308
rect 24332 10364 24396 10368
rect 24332 10308 24336 10364
rect 24336 10308 24392 10364
rect 24392 10308 24396 10364
rect 24332 10304 24396 10308
rect 24412 10364 24476 10368
rect 24412 10308 24416 10364
rect 24416 10308 24472 10364
rect 24472 10308 24476 10364
rect 24412 10304 24476 10308
rect 24492 10364 24556 10368
rect 24492 10308 24496 10364
rect 24496 10308 24552 10364
rect 24552 10308 24556 10364
rect 24492 10304 24556 10308
rect 27252 10364 27316 10368
rect 27252 10308 27256 10364
rect 27256 10308 27312 10364
rect 27312 10308 27316 10364
rect 27252 10304 27316 10308
rect 27332 10364 27396 10368
rect 27332 10308 27336 10364
rect 27336 10308 27392 10364
rect 27392 10308 27396 10364
rect 27332 10304 27396 10308
rect 27412 10364 27476 10368
rect 27412 10308 27416 10364
rect 27416 10308 27472 10364
rect 27472 10308 27476 10364
rect 27412 10304 27476 10308
rect 27492 10364 27556 10368
rect 27492 10308 27496 10364
rect 27496 10308 27552 10364
rect 27552 10308 27556 10364
rect 27492 10304 27556 10308
rect 19380 9964 19444 10028
rect 1752 9820 1816 9824
rect 1752 9764 1756 9820
rect 1756 9764 1812 9820
rect 1812 9764 1816 9820
rect 1752 9760 1816 9764
rect 1832 9820 1896 9824
rect 1832 9764 1836 9820
rect 1836 9764 1892 9820
rect 1892 9764 1896 9820
rect 1832 9760 1896 9764
rect 1912 9820 1976 9824
rect 1912 9764 1916 9820
rect 1916 9764 1972 9820
rect 1972 9764 1976 9820
rect 1912 9760 1976 9764
rect 1992 9820 2056 9824
rect 1992 9764 1996 9820
rect 1996 9764 2052 9820
rect 2052 9764 2056 9820
rect 1992 9760 2056 9764
rect 4752 9820 4816 9824
rect 4752 9764 4756 9820
rect 4756 9764 4812 9820
rect 4812 9764 4816 9820
rect 4752 9760 4816 9764
rect 4832 9820 4896 9824
rect 4832 9764 4836 9820
rect 4836 9764 4892 9820
rect 4892 9764 4896 9820
rect 4832 9760 4896 9764
rect 4912 9820 4976 9824
rect 4912 9764 4916 9820
rect 4916 9764 4972 9820
rect 4972 9764 4976 9820
rect 4912 9760 4976 9764
rect 4992 9820 5056 9824
rect 4992 9764 4996 9820
rect 4996 9764 5052 9820
rect 5052 9764 5056 9820
rect 4992 9760 5056 9764
rect 7752 9820 7816 9824
rect 7752 9764 7756 9820
rect 7756 9764 7812 9820
rect 7812 9764 7816 9820
rect 7752 9760 7816 9764
rect 7832 9820 7896 9824
rect 7832 9764 7836 9820
rect 7836 9764 7892 9820
rect 7892 9764 7896 9820
rect 7832 9760 7896 9764
rect 7912 9820 7976 9824
rect 7912 9764 7916 9820
rect 7916 9764 7972 9820
rect 7972 9764 7976 9820
rect 7912 9760 7976 9764
rect 7992 9820 8056 9824
rect 7992 9764 7996 9820
rect 7996 9764 8052 9820
rect 8052 9764 8056 9820
rect 7992 9760 8056 9764
rect 10752 9820 10816 9824
rect 10752 9764 10756 9820
rect 10756 9764 10812 9820
rect 10812 9764 10816 9820
rect 10752 9760 10816 9764
rect 10832 9820 10896 9824
rect 10832 9764 10836 9820
rect 10836 9764 10892 9820
rect 10892 9764 10896 9820
rect 10832 9760 10896 9764
rect 10912 9820 10976 9824
rect 10912 9764 10916 9820
rect 10916 9764 10972 9820
rect 10972 9764 10976 9820
rect 10912 9760 10976 9764
rect 10992 9820 11056 9824
rect 10992 9764 10996 9820
rect 10996 9764 11052 9820
rect 11052 9764 11056 9820
rect 10992 9760 11056 9764
rect 13752 9820 13816 9824
rect 13752 9764 13756 9820
rect 13756 9764 13812 9820
rect 13812 9764 13816 9820
rect 13752 9760 13816 9764
rect 13832 9820 13896 9824
rect 13832 9764 13836 9820
rect 13836 9764 13892 9820
rect 13892 9764 13896 9820
rect 13832 9760 13896 9764
rect 13912 9820 13976 9824
rect 13912 9764 13916 9820
rect 13916 9764 13972 9820
rect 13972 9764 13976 9820
rect 13912 9760 13976 9764
rect 13992 9820 14056 9824
rect 13992 9764 13996 9820
rect 13996 9764 14052 9820
rect 14052 9764 14056 9820
rect 13992 9760 14056 9764
rect 16752 9820 16816 9824
rect 16752 9764 16756 9820
rect 16756 9764 16812 9820
rect 16812 9764 16816 9820
rect 16752 9760 16816 9764
rect 16832 9820 16896 9824
rect 16832 9764 16836 9820
rect 16836 9764 16892 9820
rect 16892 9764 16896 9820
rect 16832 9760 16896 9764
rect 16912 9820 16976 9824
rect 16912 9764 16916 9820
rect 16916 9764 16972 9820
rect 16972 9764 16976 9820
rect 16912 9760 16976 9764
rect 16992 9820 17056 9824
rect 16992 9764 16996 9820
rect 16996 9764 17052 9820
rect 17052 9764 17056 9820
rect 16992 9760 17056 9764
rect 19752 9820 19816 9824
rect 19752 9764 19756 9820
rect 19756 9764 19812 9820
rect 19812 9764 19816 9820
rect 19752 9760 19816 9764
rect 19832 9820 19896 9824
rect 19832 9764 19836 9820
rect 19836 9764 19892 9820
rect 19892 9764 19896 9820
rect 19832 9760 19896 9764
rect 19912 9820 19976 9824
rect 19912 9764 19916 9820
rect 19916 9764 19972 9820
rect 19972 9764 19976 9820
rect 19912 9760 19976 9764
rect 19992 9820 20056 9824
rect 19992 9764 19996 9820
rect 19996 9764 20052 9820
rect 20052 9764 20056 9820
rect 19992 9760 20056 9764
rect 22752 9820 22816 9824
rect 22752 9764 22756 9820
rect 22756 9764 22812 9820
rect 22812 9764 22816 9820
rect 22752 9760 22816 9764
rect 22832 9820 22896 9824
rect 22832 9764 22836 9820
rect 22836 9764 22892 9820
rect 22892 9764 22896 9820
rect 22832 9760 22896 9764
rect 22912 9820 22976 9824
rect 22912 9764 22916 9820
rect 22916 9764 22972 9820
rect 22972 9764 22976 9820
rect 22912 9760 22976 9764
rect 22992 9820 23056 9824
rect 22992 9764 22996 9820
rect 22996 9764 23052 9820
rect 23052 9764 23056 9820
rect 22992 9760 23056 9764
rect 25752 9820 25816 9824
rect 25752 9764 25756 9820
rect 25756 9764 25812 9820
rect 25812 9764 25816 9820
rect 25752 9760 25816 9764
rect 25832 9820 25896 9824
rect 25832 9764 25836 9820
rect 25836 9764 25892 9820
rect 25892 9764 25896 9820
rect 25832 9760 25896 9764
rect 25912 9820 25976 9824
rect 25912 9764 25916 9820
rect 25916 9764 25972 9820
rect 25972 9764 25976 9820
rect 25912 9760 25976 9764
rect 25992 9820 26056 9824
rect 25992 9764 25996 9820
rect 25996 9764 26052 9820
rect 26052 9764 26056 9820
rect 25992 9760 26056 9764
rect 3252 9276 3316 9280
rect 3252 9220 3256 9276
rect 3256 9220 3312 9276
rect 3312 9220 3316 9276
rect 3252 9216 3316 9220
rect 3332 9276 3396 9280
rect 3332 9220 3336 9276
rect 3336 9220 3392 9276
rect 3392 9220 3396 9276
rect 3332 9216 3396 9220
rect 3412 9276 3476 9280
rect 3412 9220 3416 9276
rect 3416 9220 3472 9276
rect 3472 9220 3476 9276
rect 3412 9216 3476 9220
rect 3492 9276 3556 9280
rect 3492 9220 3496 9276
rect 3496 9220 3552 9276
rect 3552 9220 3556 9276
rect 3492 9216 3556 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 6412 9276 6476 9280
rect 6412 9220 6416 9276
rect 6416 9220 6472 9276
rect 6472 9220 6476 9276
rect 6412 9216 6476 9220
rect 6492 9276 6556 9280
rect 6492 9220 6496 9276
rect 6496 9220 6552 9276
rect 6552 9220 6556 9276
rect 6492 9216 6556 9220
rect 9252 9276 9316 9280
rect 9252 9220 9256 9276
rect 9256 9220 9312 9276
rect 9312 9220 9316 9276
rect 9252 9216 9316 9220
rect 9332 9276 9396 9280
rect 9332 9220 9336 9276
rect 9336 9220 9392 9276
rect 9392 9220 9396 9276
rect 9332 9216 9396 9220
rect 9412 9276 9476 9280
rect 9412 9220 9416 9276
rect 9416 9220 9472 9276
rect 9472 9220 9476 9276
rect 9412 9216 9476 9220
rect 9492 9276 9556 9280
rect 9492 9220 9496 9276
rect 9496 9220 9552 9276
rect 9552 9220 9556 9276
rect 9492 9216 9556 9220
rect 12252 9276 12316 9280
rect 12252 9220 12256 9276
rect 12256 9220 12312 9276
rect 12312 9220 12316 9276
rect 12252 9216 12316 9220
rect 12332 9276 12396 9280
rect 12332 9220 12336 9276
rect 12336 9220 12392 9276
rect 12392 9220 12396 9276
rect 12332 9216 12396 9220
rect 12412 9276 12476 9280
rect 12412 9220 12416 9276
rect 12416 9220 12472 9276
rect 12472 9220 12476 9276
rect 12412 9216 12476 9220
rect 12492 9276 12556 9280
rect 12492 9220 12496 9276
rect 12496 9220 12552 9276
rect 12552 9220 12556 9276
rect 12492 9216 12556 9220
rect 15252 9276 15316 9280
rect 15252 9220 15256 9276
rect 15256 9220 15312 9276
rect 15312 9220 15316 9276
rect 15252 9216 15316 9220
rect 15332 9276 15396 9280
rect 15332 9220 15336 9276
rect 15336 9220 15392 9276
rect 15392 9220 15396 9276
rect 15332 9216 15396 9220
rect 15412 9276 15476 9280
rect 15412 9220 15416 9276
rect 15416 9220 15472 9276
rect 15472 9220 15476 9276
rect 15412 9216 15476 9220
rect 15492 9276 15556 9280
rect 15492 9220 15496 9276
rect 15496 9220 15552 9276
rect 15552 9220 15556 9276
rect 15492 9216 15556 9220
rect 18252 9276 18316 9280
rect 18252 9220 18256 9276
rect 18256 9220 18312 9276
rect 18312 9220 18316 9276
rect 18252 9216 18316 9220
rect 18332 9276 18396 9280
rect 18332 9220 18336 9276
rect 18336 9220 18392 9276
rect 18392 9220 18396 9276
rect 18332 9216 18396 9220
rect 18412 9276 18476 9280
rect 18412 9220 18416 9276
rect 18416 9220 18472 9276
rect 18472 9220 18476 9276
rect 18412 9216 18476 9220
rect 18492 9276 18556 9280
rect 18492 9220 18496 9276
rect 18496 9220 18552 9276
rect 18552 9220 18556 9276
rect 18492 9216 18556 9220
rect 21252 9276 21316 9280
rect 21252 9220 21256 9276
rect 21256 9220 21312 9276
rect 21312 9220 21316 9276
rect 21252 9216 21316 9220
rect 21332 9276 21396 9280
rect 21332 9220 21336 9276
rect 21336 9220 21392 9276
rect 21392 9220 21396 9276
rect 21332 9216 21396 9220
rect 21412 9276 21476 9280
rect 21412 9220 21416 9276
rect 21416 9220 21472 9276
rect 21472 9220 21476 9276
rect 21412 9216 21476 9220
rect 21492 9276 21556 9280
rect 21492 9220 21496 9276
rect 21496 9220 21552 9276
rect 21552 9220 21556 9276
rect 21492 9216 21556 9220
rect 24252 9276 24316 9280
rect 24252 9220 24256 9276
rect 24256 9220 24312 9276
rect 24312 9220 24316 9276
rect 24252 9216 24316 9220
rect 24332 9276 24396 9280
rect 24332 9220 24336 9276
rect 24336 9220 24392 9276
rect 24392 9220 24396 9276
rect 24332 9216 24396 9220
rect 24412 9276 24476 9280
rect 24412 9220 24416 9276
rect 24416 9220 24472 9276
rect 24472 9220 24476 9276
rect 24412 9216 24476 9220
rect 24492 9276 24556 9280
rect 24492 9220 24496 9276
rect 24496 9220 24552 9276
rect 24552 9220 24556 9276
rect 24492 9216 24556 9220
rect 27252 9276 27316 9280
rect 27252 9220 27256 9276
rect 27256 9220 27312 9276
rect 27312 9220 27316 9276
rect 27252 9216 27316 9220
rect 27332 9276 27396 9280
rect 27332 9220 27336 9276
rect 27336 9220 27392 9276
rect 27392 9220 27396 9276
rect 27332 9216 27396 9220
rect 27412 9276 27476 9280
rect 27412 9220 27416 9276
rect 27416 9220 27472 9276
rect 27472 9220 27476 9276
rect 27412 9216 27476 9220
rect 27492 9276 27556 9280
rect 27492 9220 27496 9276
rect 27496 9220 27552 9276
rect 27552 9220 27556 9276
rect 27492 9216 27556 9220
rect 1752 8732 1816 8736
rect 1752 8676 1756 8732
rect 1756 8676 1812 8732
rect 1812 8676 1816 8732
rect 1752 8672 1816 8676
rect 1832 8732 1896 8736
rect 1832 8676 1836 8732
rect 1836 8676 1892 8732
rect 1892 8676 1896 8732
rect 1832 8672 1896 8676
rect 1912 8732 1976 8736
rect 1912 8676 1916 8732
rect 1916 8676 1972 8732
rect 1972 8676 1976 8732
rect 1912 8672 1976 8676
rect 1992 8732 2056 8736
rect 1992 8676 1996 8732
rect 1996 8676 2052 8732
rect 2052 8676 2056 8732
rect 1992 8672 2056 8676
rect 4752 8732 4816 8736
rect 4752 8676 4756 8732
rect 4756 8676 4812 8732
rect 4812 8676 4816 8732
rect 4752 8672 4816 8676
rect 4832 8732 4896 8736
rect 4832 8676 4836 8732
rect 4836 8676 4892 8732
rect 4892 8676 4896 8732
rect 4832 8672 4896 8676
rect 4912 8732 4976 8736
rect 4912 8676 4916 8732
rect 4916 8676 4972 8732
rect 4972 8676 4976 8732
rect 4912 8672 4976 8676
rect 4992 8732 5056 8736
rect 4992 8676 4996 8732
rect 4996 8676 5052 8732
rect 5052 8676 5056 8732
rect 4992 8672 5056 8676
rect 7752 8732 7816 8736
rect 7752 8676 7756 8732
rect 7756 8676 7812 8732
rect 7812 8676 7816 8732
rect 7752 8672 7816 8676
rect 7832 8732 7896 8736
rect 7832 8676 7836 8732
rect 7836 8676 7892 8732
rect 7892 8676 7896 8732
rect 7832 8672 7896 8676
rect 7912 8732 7976 8736
rect 7912 8676 7916 8732
rect 7916 8676 7972 8732
rect 7972 8676 7976 8732
rect 7912 8672 7976 8676
rect 7992 8732 8056 8736
rect 7992 8676 7996 8732
rect 7996 8676 8052 8732
rect 8052 8676 8056 8732
rect 7992 8672 8056 8676
rect 10752 8732 10816 8736
rect 10752 8676 10756 8732
rect 10756 8676 10812 8732
rect 10812 8676 10816 8732
rect 10752 8672 10816 8676
rect 10832 8732 10896 8736
rect 10832 8676 10836 8732
rect 10836 8676 10892 8732
rect 10892 8676 10896 8732
rect 10832 8672 10896 8676
rect 10912 8732 10976 8736
rect 10912 8676 10916 8732
rect 10916 8676 10972 8732
rect 10972 8676 10976 8732
rect 10912 8672 10976 8676
rect 10992 8732 11056 8736
rect 10992 8676 10996 8732
rect 10996 8676 11052 8732
rect 11052 8676 11056 8732
rect 10992 8672 11056 8676
rect 13752 8732 13816 8736
rect 13752 8676 13756 8732
rect 13756 8676 13812 8732
rect 13812 8676 13816 8732
rect 13752 8672 13816 8676
rect 13832 8732 13896 8736
rect 13832 8676 13836 8732
rect 13836 8676 13892 8732
rect 13892 8676 13896 8732
rect 13832 8672 13896 8676
rect 13912 8732 13976 8736
rect 13912 8676 13916 8732
rect 13916 8676 13972 8732
rect 13972 8676 13976 8732
rect 13912 8672 13976 8676
rect 13992 8732 14056 8736
rect 13992 8676 13996 8732
rect 13996 8676 14052 8732
rect 14052 8676 14056 8732
rect 13992 8672 14056 8676
rect 16752 8732 16816 8736
rect 16752 8676 16756 8732
rect 16756 8676 16812 8732
rect 16812 8676 16816 8732
rect 16752 8672 16816 8676
rect 16832 8732 16896 8736
rect 16832 8676 16836 8732
rect 16836 8676 16892 8732
rect 16892 8676 16896 8732
rect 16832 8672 16896 8676
rect 16912 8732 16976 8736
rect 16912 8676 16916 8732
rect 16916 8676 16972 8732
rect 16972 8676 16976 8732
rect 16912 8672 16976 8676
rect 16992 8732 17056 8736
rect 16992 8676 16996 8732
rect 16996 8676 17052 8732
rect 17052 8676 17056 8732
rect 16992 8672 17056 8676
rect 19752 8732 19816 8736
rect 19752 8676 19756 8732
rect 19756 8676 19812 8732
rect 19812 8676 19816 8732
rect 19752 8672 19816 8676
rect 19832 8732 19896 8736
rect 19832 8676 19836 8732
rect 19836 8676 19892 8732
rect 19892 8676 19896 8732
rect 19832 8672 19896 8676
rect 19912 8732 19976 8736
rect 19912 8676 19916 8732
rect 19916 8676 19972 8732
rect 19972 8676 19976 8732
rect 19912 8672 19976 8676
rect 19992 8732 20056 8736
rect 19992 8676 19996 8732
rect 19996 8676 20052 8732
rect 20052 8676 20056 8732
rect 19992 8672 20056 8676
rect 22752 8732 22816 8736
rect 22752 8676 22756 8732
rect 22756 8676 22812 8732
rect 22812 8676 22816 8732
rect 22752 8672 22816 8676
rect 22832 8732 22896 8736
rect 22832 8676 22836 8732
rect 22836 8676 22892 8732
rect 22892 8676 22896 8732
rect 22832 8672 22896 8676
rect 22912 8732 22976 8736
rect 22912 8676 22916 8732
rect 22916 8676 22972 8732
rect 22972 8676 22976 8732
rect 22912 8672 22976 8676
rect 22992 8732 23056 8736
rect 22992 8676 22996 8732
rect 22996 8676 23052 8732
rect 23052 8676 23056 8732
rect 22992 8672 23056 8676
rect 25752 8732 25816 8736
rect 25752 8676 25756 8732
rect 25756 8676 25812 8732
rect 25812 8676 25816 8732
rect 25752 8672 25816 8676
rect 25832 8732 25896 8736
rect 25832 8676 25836 8732
rect 25836 8676 25892 8732
rect 25892 8676 25896 8732
rect 25832 8672 25896 8676
rect 25912 8732 25976 8736
rect 25912 8676 25916 8732
rect 25916 8676 25972 8732
rect 25972 8676 25976 8732
rect 25912 8672 25976 8676
rect 25992 8732 26056 8736
rect 25992 8676 25996 8732
rect 25996 8676 26052 8732
rect 26052 8676 26056 8732
rect 25992 8672 26056 8676
rect 3252 8188 3316 8192
rect 3252 8132 3256 8188
rect 3256 8132 3312 8188
rect 3312 8132 3316 8188
rect 3252 8128 3316 8132
rect 3332 8188 3396 8192
rect 3332 8132 3336 8188
rect 3336 8132 3392 8188
rect 3392 8132 3396 8188
rect 3332 8128 3396 8132
rect 3412 8188 3476 8192
rect 3412 8132 3416 8188
rect 3416 8132 3472 8188
rect 3472 8132 3476 8188
rect 3412 8128 3476 8132
rect 3492 8188 3556 8192
rect 3492 8132 3496 8188
rect 3496 8132 3552 8188
rect 3552 8132 3556 8188
rect 3492 8128 3556 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 6412 8188 6476 8192
rect 6412 8132 6416 8188
rect 6416 8132 6472 8188
rect 6472 8132 6476 8188
rect 6412 8128 6476 8132
rect 6492 8188 6556 8192
rect 6492 8132 6496 8188
rect 6496 8132 6552 8188
rect 6552 8132 6556 8188
rect 6492 8128 6556 8132
rect 9252 8188 9316 8192
rect 9252 8132 9256 8188
rect 9256 8132 9312 8188
rect 9312 8132 9316 8188
rect 9252 8128 9316 8132
rect 9332 8188 9396 8192
rect 9332 8132 9336 8188
rect 9336 8132 9392 8188
rect 9392 8132 9396 8188
rect 9332 8128 9396 8132
rect 9412 8188 9476 8192
rect 9412 8132 9416 8188
rect 9416 8132 9472 8188
rect 9472 8132 9476 8188
rect 9412 8128 9476 8132
rect 9492 8188 9556 8192
rect 9492 8132 9496 8188
rect 9496 8132 9552 8188
rect 9552 8132 9556 8188
rect 9492 8128 9556 8132
rect 12252 8188 12316 8192
rect 12252 8132 12256 8188
rect 12256 8132 12312 8188
rect 12312 8132 12316 8188
rect 12252 8128 12316 8132
rect 12332 8188 12396 8192
rect 12332 8132 12336 8188
rect 12336 8132 12392 8188
rect 12392 8132 12396 8188
rect 12332 8128 12396 8132
rect 12412 8188 12476 8192
rect 12412 8132 12416 8188
rect 12416 8132 12472 8188
rect 12472 8132 12476 8188
rect 12412 8128 12476 8132
rect 12492 8188 12556 8192
rect 12492 8132 12496 8188
rect 12496 8132 12552 8188
rect 12552 8132 12556 8188
rect 12492 8128 12556 8132
rect 15252 8188 15316 8192
rect 15252 8132 15256 8188
rect 15256 8132 15312 8188
rect 15312 8132 15316 8188
rect 15252 8128 15316 8132
rect 15332 8188 15396 8192
rect 15332 8132 15336 8188
rect 15336 8132 15392 8188
rect 15392 8132 15396 8188
rect 15332 8128 15396 8132
rect 15412 8188 15476 8192
rect 15412 8132 15416 8188
rect 15416 8132 15472 8188
rect 15472 8132 15476 8188
rect 15412 8128 15476 8132
rect 15492 8188 15556 8192
rect 15492 8132 15496 8188
rect 15496 8132 15552 8188
rect 15552 8132 15556 8188
rect 15492 8128 15556 8132
rect 18252 8188 18316 8192
rect 18252 8132 18256 8188
rect 18256 8132 18312 8188
rect 18312 8132 18316 8188
rect 18252 8128 18316 8132
rect 18332 8188 18396 8192
rect 18332 8132 18336 8188
rect 18336 8132 18392 8188
rect 18392 8132 18396 8188
rect 18332 8128 18396 8132
rect 18412 8188 18476 8192
rect 18412 8132 18416 8188
rect 18416 8132 18472 8188
rect 18472 8132 18476 8188
rect 18412 8128 18476 8132
rect 18492 8188 18556 8192
rect 18492 8132 18496 8188
rect 18496 8132 18552 8188
rect 18552 8132 18556 8188
rect 18492 8128 18556 8132
rect 21252 8188 21316 8192
rect 21252 8132 21256 8188
rect 21256 8132 21312 8188
rect 21312 8132 21316 8188
rect 21252 8128 21316 8132
rect 21332 8188 21396 8192
rect 21332 8132 21336 8188
rect 21336 8132 21392 8188
rect 21392 8132 21396 8188
rect 21332 8128 21396 8132
rect 21412 8188 21476 8192
rect 21412 8132 21416 8188
rect 21416 8132 21472 8188
rect 21472 8132 21476 8188
rect 21412 8128 21476 8132
rect 21492 8188 21556 8192
rect 21492 8132 21496 8188
rect 21496 8132 21552 8188
rect 21552 8132 21556 8188
rect 21492 8128 21556 8132
rect 24252 8188 24316 8192
rect 24252 8132 24256 8188
rect 24256 8132 24312 8188
rect 24312 8132 24316 8188
rect 24252 8128 24316 8132
rect 24332 8188 24396 8192
rect 24332 8132 24336 8188
rect 24336 8132 24392 8188
rect 24392 8132 24396 8188
rect 24332 8128 24396 8132
rect 24412 8188 24476 8192
rect 24412 8132 24416 8188
rect 24416 8132 24472 8188
rect 24472 8132 24476 8188
rect 24412 8128 24476 8132
rect 24492 8188 24556 8192
rect 24492 8132 24496 8188
rect 24496 8132 24552 8188
rect 24552 8132 24556 8188
rect 24492 8128 24556 8132
rect 27252 8188 27316 8192
rect 27252 8132 27256 8188
rect 27256 8132 27312 8188
rect 27312 8132 27316 8188
rect 27252 8128 27316 8132
rect 27332 8188 27396 8192
rect 27332 8132 27336 8188
rect 27336 8132 27392 8188
rect 27392 8132 27396 8188
rect 27332 8128 27396 8132
rect 27412 8188 27476 8192
rect 27412 8132 27416 8188
rect 27416 8132 27472 8188
rect 27472 8132 27476 8188
rect 27412 8128 27476 8132
rect 27492 8188 27556 8192
rect 27492 8132 27496 8188
rect 27496 8132 27552 8188
rect 27552 8132 27556 8188
rect 27492 8128 27556 8132
rect 1752 7644 1816 7648
rect 1752 7588 1756 7644
rect 1756 7588 1812 7644
rect 1812 7588 1816 7644
rect 1752 7584 1816 7588
rect 1832 7644 1896 7648
rect 1832 7588 1836 7644
rect 1836 7588 1892 7644
rect 1892 7588 1896 7644
rect 1832 7584 1896 7588
rect 1912 7644 1976 7648
rect 1912 7588 1916 7644
rect 1916 7588 1972 7644
rect 1972 7588 1976 7644
rect 1912 7584 1976 7588
rect 1992 7644 2056 7648
rect 1992 7588 1996 7644
rect 1996 7588 2052 7644
rect 2052 7588 2056 7644
rect 1992 7584 2056 7588
rect 4752 7644 4816 7648
rect 4752 7588 4756 7644
rect 4756 7588 4812 7644
rect 4812 7588 4816 7644
rect 4752 7584 4816 7588
rect 4832 7644 4896 7648
rect 4832 7588 4836 7644
rect 4836 7588 4892 7644
rect 4892 7588 4896 7644
rect 4832 7584 4896 7588
rect 4912 7644 4976 7648
rect 4912 7588 4916 7644
rect 4916 7588 4972 7644
rect 4972 7588 4976 7644
rect 4912 7584 4976 7588
rect 4992 7644 5056 7648
rect 4992 7588 4996 7644
rect 4996 7588 5052 7644
rect 5052 7588 5056 7644
rect 4992 7584 5056 7588
rect 7752 7644 7816 7648
rect 7752 7588 7756 7644
rect 7756 7588 7812 7644
rect 7812 7588 7816 7644
rect 7752 7584 7816 7588
rect 7832 7644 7896 7648
rect 7832 7588 7836 7644
rect 7836 7588 7892 7644
rect 7892 7588 7896 7644
rect 7832 7584 7896 7588
rect 7912 7644 7976 7648
rect 7912 7588 7916 7644
rect 7916 7588 7972 7644
rect 7972 7588 7976 7644
rect 7912 7584 7976 7588
rect 7992 7644 8056 7648
rect 7992 7588 7996 7644
rect 7996 7588 8052 7644
rect 8052 7588 8056 7644
rect 7992 7584 8056 7588
rect 10752 7644 10816 7648
rect 10752 7588 10756 7644
rect 10756 7588 10812 7644
rect 10812 7588 10816 7644
rect 10752 7584 10816 7588
rect 10832 7644 10896 7648
rect 10832 7588 10836 7644
rect 10836 7588 10892 7644
rect 10892 7588 10896 7644
rect 10832 7584 10896 7588
rect 10912 7644 10976 7648
rect 10912 7588 10916 7644
rect 10916 7588 10972 7644
rect 10972 7588 10976 7644
rect 10912 7584 10976 7588
rect 10992 7644 11056 7648
rect 10992 7588 10996 7644
rect 10996 7588 11052 7644
rect 11052 7588 11056 7644
rect 10992 7584 11056 7588
rect 13752 7644 13816 7648
rect 13752 7588 13756 7644
rect 13756 7588 13812 7644
rect 13812 7588 13816 7644
rect 13752 7584 13816 7588
rect 13832 7644 13896 7648
rect 13832 7588 13836 7644
rect 13836 7588 13892 7644
rect 13892 7588 13896 7644
rect 13832 7584 13896 7588
rect 13912 7644 13976 7648
rect 13912 7588 13916 7644
rect 13916 7588 13972 7644
rect 13972 7588 13976 7644
rect 13912 7584 13976 7588
rect 13992 7644 14056 7648
rect 13992 7588 13996 7644
rect 13996 7588 14052 7644
rect 14052 7588 14056 7644
rect 13992 7584 14056 7588
rect 16752 7644 16816 7648
rect 16752 7588 16756 7644
rect 16756 7588 16812 7644
rect 16812 7588 16816 7644
rect 16752 7584 16816 7588
rect 16832 7644 16896 7648
rect 16832 7588 16836 7644
rect 16836 7588 16892 7644
rect 16892 7588 16896 7644
rect 16832 7584 16896 7588
rect 16912 7644 16976 7648
rect 16912 7588 16916 7644
rect 16916 7588 16972 7644
rect 16972 7588 16976 7644
rect 16912 7584 16976 7588
rect 16992 7644 17056 7648
rect 16992 7588 16996 7644
rect 16996 7588 17052 7644
rect 17052 7588 17056 7644
rect 16992 7584 17056 7588
rect 19752 7644 19816 7648
rect 19752 7588 19756 7644
rect 19756 7588 19812 7644
rect 19812 7588 19816 7644
rect 19752 7584 19816 7588
rect 19832 7644 19896 7648
rect 19832 7588 19836 7644
rect 19836 7588 19892 7644
rect 19892 7588 19896 7644
rect 19832 7584 19896 7588
rect 19912 7644 19976 7648
rect 19912 7588 19916 7644
rect 19916 7588 19972 7644
rect 19972 7588 19976 7644
rect 19912 7584 19976 7588
rect 19992 7644 20056 7648
rect 19992 7588 19996 7644
rect 19996 7588 20052 7644
rect 20052 7588 20056 7644
rect 19992 7584 20056 7588
rect 22752 7644 22816 7648
rect 22752 7588 22756 7644
rect 22756 7588 22812 7644
rect 22812 7588 22816 7644
rect 22752 7584 22816 7588
rect 22832 7644 22896 7648
rect 22832 7588 22836 7644
rect 22836 7588 22892 7644
rect 22892 7588 22896 7644
rect 22832 7584 22896 7588
rect 22912 7644 22976 7648
rect 22912 7588 22916 7644
rect 22916 7588 22972 7644
rect 22972 7588 22976 7644
rect 22912 7584 22976 7588
rect 22992 7644 23056 7648
rect 22992 7588 22996 7644
rect 22996 7588 23052 7644
rect 23052 7588 23056 7644
rect 22992 7584 23056 7588
rect 25752 7644 25816 7648
rect 25752 7588 25756 7644
rect 25756 7588 25812 7644
rect 25812 7588 25816 7644
rect 25752 7584 25816 7588
rect 25832 7644 25896 7648
rect 25832 7588 25836 7644
rect 25836 7588 25892 7644
rect 25892 7588 25896 7644
rect 25832 7584 25896 7588
rect 25912 7644 25976 7648
rect 25912 7588 25916 7644
rect 25916 7588 25972 7644
rect 25972 7588 25976 7644
rect 25912 7584 25976 7588
rect 25992 7644 26056 7648
rect 25992 7588 25996 7644
rect 25996 7588 26052 7644
rect 26052 7588 26056 7644
rect 25992 7584 26056 7588
rect 3252 7100 3316 7104
rect 3252 7044 3256 7100
rect 3256 7044 3312 7100
rect 3312 7044 3316 7100
rect 3252 7040 3316 7044
rect 3332 7100 3396 7104
rect 3332 7044 3336 7100
rect 3336 7044 3392 7100
rect 3392 7044 3396 7100
rect 3332 7040 3396 7044
rect 3412 7100 3476 7104
rect 3412 7044 3416 7100
rect 3416 7044 3472 7100
rect 3472 7044 3476 7100
rect 3412 7040 3476 7044
rect 3492 7100 3556 7104
rect 3492 7044 3496 7100
rect 3496 7044 3552 7100
rect 3552 7044 3556 7100
rect 3492 7040 3556 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 6412 7100 6476 7104
rect 6412 7044 6416 7100
rect 6416 7044 6472 7100
rect 6472 7044 6476 7100
rect 6412 7040 6476 7044
rect 6492 7100 6556 7104
rect 6492 7044 6496 7100
rect 6496 7044 6552 7100
rect 6552 7044 6556 7100
rect 6492 7040 6556 7044
rect 9252 7100 9316 7104
rect 9252 7044 9256 7100
rect 9256 7044 9312 7100
rect 9312 7044 9316 7100
rect 9252 7040 9316 7044
rect 9332 7100 9396 7104
rect 9332 7044 9336 7100
rect 9336 7044 9392 7100
rect 9392 7044 9396 7100
rect 9332 7040 9396 7044
rect 9412 7100 9476 7104
rect 9412 7044 9416 7100
rect 9416 7044 9472 7100
rect 9472 7044 9476 7100
rect 9412 7040 9476 7044
rect 9492 7100 9556 7104
rect 9492 7044 9496 7100
rect 9496 7044 9552 7100
rect 9552 7044 9556 7100
rect 9492 7040 9556 7044
rect 12252 7100 12316 7104
rect 12252 7044 12256 7100
rect 12256 7044 12312 7100
rect 12312 7044 12316 7100
rect 12252 7040 12316 7044
rect 12332 7100 12396 7104
rect 12332 7044 12336 7100
rect 12336 7044 12392 7100
rect 12392 7044 12396 7100
rect 12332 7040 12396 7044
rect 12412 7100 12476 7104
rect 12412 7044 12416 7100
rect 12416 7044 12472 7100
rect 12472 7044 12476 7100
rect 12412 7040 12476 7044
rect 12492 7100 12556 7104
rect 12492 7044 12496 7100
rect 12496 7044 12552 7100
rect 12552 7044 12556 7100
rect 12492 7040 12556 7044
rect 15252 7100 15316 7104
rect 15252 7044 15256 7100
rect 15256 7044 15312 7100
rect 15312 7044 15316 7100
rect 15252 7040 15316 7044
rect 15332 7100 15396 7104
rect 15332 7044 15336 7100
rect 15336 7044 15392 7100
rect 15392 7044 15396 7100
rect 15332 7040 15396 7044
rect 15412 7100 15476 7104
rect 15412 7044 15416 7100
rect 15416 7044 15472 7100
rect 15472 7044 15476 7100
rect 15412 7040 15476 7044
rect 15492 7100 15556 7104
rect 15492 7044 15496 7100
rect 15496 7044 15552 7100
rect 15552 7044 15556 7100
rect 15492 7040 15556 7044
rect 18252 7100 18316 7104
rect 18252 7044 18256 7100
rect 18256 7044 18312 7100
rect 18312 7044 18316 7100
rect 18252 7040 18316 7044
rect 18332 7100 18396 7104
rect 18332 7044 18336 7100
rect 18336 7044 18392 7100
rect 18392 7044 18396 7100
rect 18332 7040 18396 7044
rect 18412 7100 18476 7104
rect 18412 7044 18416 7100
rect 18416 7044 18472 7100
rect 18472 7044 18476 7100
rect 18412 7040 18476 7044
rect 18492 7100 18556 7104
rect 18492 7044 18496 7100
rect 18496 7044 18552 7100
rect 18552 7044 18556 7100
rect 18492 7040 18556 7044
rect 21252 7100 21316 7104
rect 21252 7044 21256 7100
rect 21256 7044 21312 7100
rect 21312 7044 21316 7100
rect 21252 7040 21316 7044
rect 21332 7100 21396 7104
rect 21332 7044 21336 7100
rect 21336 7044 21392 7100
rect 21392 7044 21396 7100
rect 21332 7040 21396 7044
rect 21412 7100 21476 7104
rect 21412 7044 21416 7100
rect 21416 7044 21472 7100
rect 21472 7044 21476 7100
rect 21412 7040 21476 7044
rect 21492 7100 21556 7104
rect 21492 7044 21496 7100
rect 21496 7044 21552 7100
rect 21552 7044 21556 7100
rect 21492 7040 21556 7044
rect 24252 7100 24316 7104
rect 24252 7044 24256 7100
rect 24256 7044 24312 7100
rect 24312 7044 24316 7100
rect 24252 7040 24316 7044
rect 24332 7100 24396 7104
rect 24332 7044 24336 7100
rect 24336 7044 24392 7100
rect 24392 7044 24396 7100
rect 24332 7040 24396 7044
rect 24412 7100 24476 7104
rect 24412 7044 24416 7100
rect 24416 7044 24472 7100
rect 24472 7044 24476 7100
rect 24412 7040 24476 7044
rect 24492 7100 24556 7104
rect 24492 7044 24496 7100
rect 24496 7044 24552 7100
rect 24552 7044 24556 7100
rect 24492 7040 24556 7044
rect 27252 7100 27316 7104
rect 27252 7044 27256 7100
rect 27256 7044 27312 7100
rect 27312 7044 27316 7100
rect 27252 7040 27316 7044
rect 27332 7100 27396 7104
rect 27332 7044 27336 7100
rect 27336 7044 27392 7100
rect 27392 7044 27396 7100
rect 27332 7040 27396 7044
rect 27412 7100 27476 7104
rect 27412 7044 27416 7100
rect 27416 7044 27472 7100
rect 27472 7044 27476 7100
rect 27412 7040 27476 7044
rect 27492 7100 27556 7104
rect 27492 7044 27496 7100
rect 27496 7044 27552 7100
rect 27552 7044 27556 7100
rect 27492 7040 27556 7044
rect 1752 6556 1816 6560
rect 1752 6500 1756 6556
rect 1756 6500 1812 6556
rect 1812 6500 1816 6556
rect 1752 6496 1816 6500
rect 1832 6556 1896 6560
rect 1832 6500 1836 6556
rect 1836 6500 1892 6556
rect 1892 6500 1896 6556
rect 1832 6496 1896 6500
rect 1912 6556 1976 6560
rect 1912 6500 1916 6556
rect 1916 6500 1972 6556
rect 1972 6500 1976 6556
rect 1912 6496 1976 6500
rect 1992 6556 2056 6560
rect 1992 6500 1996 6556
rect 1996 6500 2052 6556
rect 2052 6500 2056 6556
rect 1992 6496 2056 6500
rect 4752 6556 4816 6560
rect 4752 6500 4756 6556
rect 4756 6500 4812 6556
rect 4812 6500 4816 6556
rect 4752 6496 4816 6500
rect 4832 6556 4896 6560
rect 4832 6500 4836 6556
rect 4836 6500 4892 6556
rect 4892 6500 4896 6556
rect 4832 6496 4896 6500
rect 4912 6556 4976 6560
rect 4912 6500 4916 6556
rect 4916 6500 4972 6556
rect 4972 6500 4976 6556
rect 4912 6496 4976 6500
rect 4992 6556 5056 6560
rect 4992 6500 4996 6556
rect 4996 6500 5052 6556
rect 5052 6500 5056 6556
rect 4992 6496 5056 6500
rect 7752 6556 7816 6560
rect 7752 6500 7756 6556
rect 7756 6500 7812 6556
rect 7812 6500 7816 6556
rect 7752 6496 7816 6500
rect 7832 6556 7896 6560
rect 7832 6500 7836 6556
rect 7836 6500 7892 6556
rect 7892 6500 7896 6556
rect 7832 6496 7896 6500
rect 7912 6556 7976 6560
rect 7912 6500 7916 6556
rect 7916 6500 7972 6556
rect 7972 6500 7976 6556
rect 7912 6496 7976 6500
rect 7992 6556 8056 6560
rect 7992 6500 7996 6556
rect 7996 6500 8052 6556
rect 8052 6500 8056 6556
rect 7992 6496 8056 6500
rect 10752 6556 10816 6560
rect 10752 6500 10756 6556
rect 10756 6500 10812 6556
rect 10812 6500 10816 6556
rect 10752 6496 10816 6500
rect 10832 6556 10896 6560
rect 10832 6500 10836 6556
rect 10836 6500 10892 6556
rect 10892 6500 10896 6556
rect 10832 6496 10896 6500
rect 10912 6556 10976 6560
rect 10912 6500 10916 6556
rect 10916 6500 10972 6556
rect 10972 6500 10976 6556
rect 10912 6496 10976 6500
rect 10992 6556 11056 6560
rect 10992 6500 10996 6556
rect 10996 6500 11052 6556
rect 11052 6500 11056 6556
rect 10992 6496 11056 6500
rect 13752 6556 13816 6560
rect 13752 6500 13756 6556
rect 13756 6500 13812 6556
rect 13812 6500 13816 6556
rect 13752 6496 13816 6500
rect 13832 6556 13896 6560
rect 13832 6500 13836 6556
rect 13836 6500 13892 6556
rect 13892 6500 13896 6556
rect 13832 6496 13896 6500
rect 13912 6556 13976 6560
rect 13912 6500 13916 6556
rect 13916 6500 13972 6556
rect 13972 6500 13976 6556
rect 13912 6496 13976 6500
rect 13992 6556 14056 6560
rect 13992 6500 13996 6556
rect 13996 6500 14052 6556
rect 14052 6500 14056 6556
rect 13992 6496 14056 6500
rect 16752 6556 16816 6560
rect 16752 6500 16756 6556
rect 16756 6500 16812 6556
rect 16812 6500 16816 6556
rect 16752 6496 16816 6500
rect 16832 6556 16896 6560
rect 16832 6500 16836 6556
rect 16836 6500 16892 6556
rect 16892 6500 16896 6556
rect 16832 6496 16896 6500
rect 16912 6556 16976 6560
rect 16912 6500 16916 6556
rect 16916 6500 16972 6556
rect 16972 6500 16976 6556
rect 16912 6496 16976 6500
rect 16992 6556 17056 6560
rect 16992 6500 16996 6556
rect 16996 6500 17052 6556
rect 17052 6500 17056 6556
rect 16992 6496 17056 6500
rect 19752 6556 19816 6560
rect 19752 6500 19756 6556
rect 19756 6500 19812 6556
rect 19812 6500 19816 6556
rect 19752 6496 19816 6500
rect 19832 6556 19896 6560
rect 19832 6500 19836 6556
rect 19836 6500 19892 6556
rect 19892 6500 19896 6556
rect 19832 6496 19896 6500
rect 19912 6556 19976 6560
rect 19912 6500 19916 6556
rect 19916 6500 19972 6556
rect 19972 6500 19976 6556
rect 19912 6496 19976 6500
rect 19992 6556 20056 6560
rect 19992 6500 19996 6556
rect 19996 6500 20052 6556
rect 20052 6500 20056 6556
rect 19992 6496 20056 6500
rect 22752 6556 22816 6560
rect 22752 6500 22756 6556
rect 22756 6500 22812 6556
rect 22812 6500 22816 6556
rect 22752 6496 22816 6500
rect 22832 6556 22896 6560
rect 22832 6500 22836 6556
rect 22836 6500 22892 6556
rect 22892 6500 22896 6556
rect 22832 6496 22896 6500
rect 22912 6556 22976 6560
rect 22912 6500 22916 6556
rect 22916 6500 22972 6556
rect 22972 6500 22976 6556
rect 22912 6496 22976 6500
rect 22992 6556 23056 6560
rect 22992 6500 22996 6556
rect 22996 6500 23052 6556
rect 23052 6500 23056 6556
rect 22992 6496 23056 6500
rect 25752 6556 25816 6560
rect 25752 6500 25756 6556
rect 25756 6500 25812 6556
rect 25812 6500 25816 6556
rect 25752 6496 25816 6500
rect 25832 6556 25896 6560
rect 25832 6500 25836 6556
rect 25836 6500 25892 6556
rect 25892 6500 25896 6556
rect 25832 6496 25896 6500
rect 25912 6556 25976 6560
rect 25912 6500 25916 6556
rect 25916 6500 25972 6556
rect 25972 6500 25976 6556
rect 25912 6496 25976 6500
rect 25992 6556 26056 6560
rect 25992 6500 25996 6556
rect 25996 6500 26052 6556
rect 26052 6500 26056 6556
rect 25992 6496 26056 6500
rect 3252 6012 3316 6016
rect 3252 5956 3256 6012
rect 3256 5956 3312 6012
rect 3312 5956 3316 6012
rect 3252 5952 3316 5956
rect 3332 6012 3396 6016
rect 3332 5956 3336 6012
rect 3336 5956 3392 6012
rect 3392 5956 3396 6012
rect 3332 5952 3396 5956
rect 3412 6012 3476 6016
rect 3412 5956 3416 6012
rect 3416 5956 3472 6012
rect 3472 5956 3476 6012
rect 3412 5952 3476 5956
rect 3492 6012 3556 6016
rect 3492 5956 3496 6012
rect 3496 5956 3552 6012
rect 3552 5956 3556 6012
rect 3492 5952 3556 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 6412 6012 6476 6016
rect 6412 5956 6416 6012
rect 6416 5956 6472 6012
rect 6472 5956 6476 6012
rect 6412 5952 6476 5956
rect 6492 6012 6556 6016
rect 6492 5956 6496 6012
rect 6496 5956 6552 6012
rect 6552 5956 6556 6012
rect 6492 5952 6556 5956
rect 9252 6012 9316 6016
rect 9252 5956 9256 6012
rect 9256 5956 9312 6012
rect 9312 5956 9316 6012
rect 9252 5952 9316 5956
rect 9332 6012 9396 6016
rect 9332 5956 9336 6012
rect 9336 5956 9392 6012
rect 9392 5956 9396 6012
rect 9332 5952 9396 5956
rect 9412 6012 9476 6016
rect 9412 5956 9416 6012
rect 9416 5956 9472 6012
rect 9472 5956 9476 6012
rect 9412 5952 9476 5956
rect 9492 6012 9556 6016
rect 9492 5956 9496 6012
rect 9496 5956 9552 6012
rect 9552 5956 9556 6012
rect 9492 5952 9556 5956
rect 12252 6012 12316 6016
rect 12252 5956 12256 6012
rect 12256 5956 12312 6012
rect 12312 5956 12316 6012
rect 12252 5952 12316 5956
rect 12332 6012 12396 6016
rect 12332 5956 12336 6012
rect 12336 5956 12392 6012
rect 12392 5956 12396 6012
rect 12332 5952 12396 5956
rect 12412 6012 12476 6016
rect 12412 5956 12416 6012
rect 12416 5956 12472 6012
rect 12472 5956 12476 6012
rect 12412 5952 12476 5956
rect 12492 6012 12556 6016
rect 12492 5956 12496 6012
rect 12496 5956 12552 6012
rect 12552 5956 12556 6012
rect 12492 5952 12556 5956
rect 15252 6012 15316 6016
rect 15252 5956 15256 6012
rect 15256 5956 15312 6012
rect 15312 5956 15316 6012
rect 15252 5952 15316 5956
rect 15332 6012 15396 6016
rect 15332 5956 15336 6012
rect 15336 5956 15392 6012
rect 15392 5956 15396 6012
rect 15332 5952 15396 5956
rect 15412 6012 15476 6016
rect 15412 5956 15416 6012
rect 15416 5956 15472 6012
rect 15472 5956 15476 6012
rect 15412 5952 15476 5956
rect 15492 6012 15556 6016
rect 15492 5956 15496 6012
rect 15496 5956 15552 6012
rect 15552 5956 15556 6012
rect 15492 5952 15556 5956
rect 18252 6012 18316 6016
rect 18252 5956 18256 6012
rect 18256 5956 18312 6012
rect 18312 5956 18316 6012
rect 18252 5952 18316 5956
rect 18332 6012 18396 6016
rect 18332 5956 18336 6012
rect 18336 5956 18392 6012
rect 18392 5956 18396 6012
rect 18332 5952 18396 5956
rect 18412 6012 18476 6016
rect 18412 5956 18416 6012
rect 18416 5956 18472 6012
rect 18472 5956 18476 6012
rect 18412 5952 18476 5956
rect 18492 6012 18556 6016
rect 18492 5956 18496 6012
rect 18496 5956 18552 6012
rect 18552 5956 18556 6012
rect 18492 5952 18556 5956
rect 21252 6012 21316 6016
rect 21252 5956 21256 6012
rect 21256 5956 21312 6012
rect 21312 5956 21316 6012
rect 21252 5952 21316 5956
rect 21332 6012 21396 6016
rect 21332 5956 21336 6012
rect 21336 5956 21392 6012
rect 21392 5956 21396 6012
rect 21332 5952 21396 5956
rect 21412 6012 21476 6016
rect 21412 5956 21416 6012
rect 21416 5956 21472 6012
rect 21472 5956 21476 6012
rect 21412 5952 21476 5956
rect 21492 6012 21556 6016
rect 21492 5956 21496 6012
rect 21496 5956 21552 6012
rect 21552 5956 21556 6012
rect 21492 5952 21556 5956
rect 24252 6012 24316 6016
rect 24252 5956 24256 6012
rect 24256 5956 24312 6012
rect 24312 5956 24316 6012
rect 24252 5952 24316 5956
rect 24332 6012 24396 6016
rect 24332 5956 24336 6012
rect 24336 5956 24392 6012
rect 24392 5956 24396 6012
rect 24332 5952 24396 5956
rect 24412 6012 24476 6016
rect 24412 5956 24416 6012
rect 24416 5956 24472 6012
rect 24472 5956 24476 6012
rect 24412 5952 24476 5956
rect 24492 6012 24556 6016
rect 24492 5956 24496 6012
rect 24496 5956 24552 6012
rect 24552 5956 24556 6012
rect 24492 5952 24556 5956
rect 27252 6012 27316 6016
rect 27252 5956 27256 6012
rect 27256 5956 27312 6012
rect 27312 5956 27316 6012
rect 27252 5952 27316 5956
rect 27332 6012 27396 6016
rect 27332 5956 27336 6012
rect 27336 5956 27392 6012
rect 27392 5956 27396 6012
rect 27332 5952 27396 5956
rect 27412 6012 27476 6016
rect 27412 5956 27416 6012
rect 27416 5956 27472 6012
rect 27472 5956 27476 6012
rect 27412 5952 27476 5956
rect 27492 6012 27556 6016
rect 27492 5956 27496 6012
rect 27496 5956 27552 6012
rect 27552 5956 27556 6012
rect 27492 5952 27556 5956
rect 1752 5468 1816 5472
rect 1752 5412 1756 5468
rect 1756 5412 1812 5468
rect 1812 5412 1816 5468
rect 1752 5408 1816 5412
rect 1832 5468 1896 5472
rect 1832 5412 1836 5468
rect 1836 5412 1892 5468
rect 1892 5412 1896 5468
rect 1832 5408 1896 5412
rect 1912 5468 1976 5472
rect 1912 5412 1916 5468
rect 1916 5412 1972 5468
rect 1972 5412 1976 5468
rect 1912 5408 1976 5412
rect 1992 5468 2056 5472
rect 1992 5412 1996 5468
rect 1996 5412 2052 5468
rect 2052 5412 2056 5468
rect 1992 5408 2056 5412
rect 4752 5468 4816 5472
rect 4752 5412 4756 5468
rect 4756 5412 4812 5468
rect 4812 5412 4816 5468
rect 4752 5408 4816 5412
rect 4832 5468 4896 5472
rect 4832 5412 4836 5468
rect 4836 5412 4892 5468
rect 4892 5412 4896 5468
rect 4832 5408 4896 5412
rect 4912 5468 4976 5472
rect 4912 5412 4916 5468
rect 4916 5412 4972 5468
rect 4972 5412 4976 5468
rect 4912 5408 4976 5412
rect 4992 5468 5056 5472
rect 4992 5412 4996 5468
rect 4996 5412 5052 5468
rect 5052 5412 5056 5468
rect 4992 5408 5056 5412
rect 7752 5468 7816 5472
rect 7752 5412 7756 5468
rect 7756 5412 7812 5468
rect 7812 5412 7816 5468
rect 7752 5408 7816 5412
rect 7832 5468 7896 5472
rect 7832 5412 7836 5468
rect 7836 5412 7892 5468
rect 7892 5412 7896 5468
rect 7832 5408 7896 5412
rect 7912 5468 7976 5472
rect 7912 5412 7916 5468
rect 7916 5412 7972 5468
rect 7972 5412 7976 5468
rect 7912 5408 7976 5412
rect 7992 5468 8056 5472
rect 7992 5412 7996 5468
rect 7996 5412 8052 5468
rect 8052 5412 8056 5468
rect 7992 5408 8056 5412
rect 10752 5468 10816 5472
rect 10752 5412 10756 5468
rect 10756 5412 10812 5468
rect 10812 5412 10816 5468
rect 10752 5408 10816 5412
rect 10832 5468 10896 5472
rect 10832 5412 10836 5468
rect 10836 5412 10892 5468
rect 10892 5412 10896 5468
rect 10832 5408 10896 5412
rect 10912 5468 10976 5472
rect 10912 5412 10916 5468
rect 10916 5412 10972 5468
rect 10972 5412 10976 5468
rect 10912 5408 10976 5412
rect 10992 5468 11056 5472
rect 10992 5412 10996 5468
rect 10996 5412 11052 5468
rect 11052 5412 11056 5468
rect 10992 5408 11056 5412
rect 13752 5468 13816 5472
rect 13752 5412 13756 5468
rect 13756 5412 13812 5468
rect 13812 5412 13816 5468
rect 13752 5408 13816 5412
rect 13832 5468 13896 5472
rect 13832 5412 13836 5468
rect 13836 5412 13892 5468
rect 13892 5412 13896 5468
rect 13832 5408 13896 5412
rect 13912 5468 13976 5472
rect 13912 5412 13916 5468
rect 13916 5412 13972 5468
rect 13972 5412 13976 5468
rect 13912 5408 13976 5412
rect 13992 5468 14056 5472
rect 13992 5412 13996 5468
rect 13996 5412 14052 5468
rect 14052 5412 14056 5468
rect 13992 5408 14056 5412
rect 16752 5468 16816 5472
rect 16752 5412 16756 5468
rect 16756 5412 16812 5468
rect 16812 5412 16816 5468
rect 16752 5408 16816 5412
rect 16832 5468 16896 5472
rect 16832 5412 16836 5468
rect 16836 5412 16892 5468
rect 16892 5412 16896 5468
rect 16832 5408 16896 5412
rect 16912 5468 16976 5472
rect 16912 5412 16916 5468
rect 16916 5412 16972 5468
rect 16972 5412 16976 5468
rect 16912 5408 16976 5412
rect 16992 5468 17056 5472
rect 16992 5412 16996 5468
rect 16996 5412 17052 5468
rect 17052 5412 17056 5468
rect 16992 5408 17056 5412
rect 19752 5468 19816 5472
rect 19752 5412 19756 5468
rect 19756 5412 19812 5468
rect 19812 5412 19816 5468
rect 19752 5408 19816 5412
rect 19832 5468 19896 5472
rect 19832 5412 19836 5468
rect 19836 5412 19892 5468
rect 19892 5412 19896 5468
rect 19832 5408 19896 5412
rect 19912 5468 19976 5472
rect 19912 5412 19916 5468
rect 19916 5412 19972 5468
rect 19972 5412 19976 5468
rect 19912 5408 19976 5412
rect 19992 5468 20056 5472
rect 19992 5412 19996 5468
rect 19996 5412 20052 5468
rect 20052 5412 20056 5468
rect 19992 5408 20056 5412
rect 22752 5468 22816 5472
rect 22752 5412 22756 5468
rect 22756 5412 22812 5468
rect 22812 5412 22816 5468
rect 22752 5408 22816 5412
rect 22832 5468 22896 5472
rect 22832 5412 22836 5468
rect 22836 5412 22892 5468
rect 22892 5412 22896 5468
rect 22832 5408 22896 5412
rect 22912 5468 22976 5472
rect 22912 5412 22916 5468
rect 22916 5412 22972 5468
rect 22972 5412 22976 5468
rect 22912 5408 22976 5412
rect 22992 5468 23056 5472
rect 22992 5412 22996 5468
rect 22996 5412 23052 5468
rect 23052 5412 23056 5468
rect 22992 5408 23056 5412
rect 25752 5468 25816 5472
rect 25752 5412 25756 5468
rect 25756 5412 25812 5468
rect 25812 5412 25816 5468
rect 25752 5408 25816 5412
rect 25832 5468 25896 5472
rect 25832 5412 25836 5468
rect 25836 5412 25892 5468
rect 25892 5412 25896 5468
rect 25832 5408 25896 5412
rect 25912 5468 25976 5472
rect 25912 5412 25916 5468
rect 25916 5412 25972 5468
rect 25972 5412 25976 5468
rect 25912 5408 25976 5412
rect 25992 5468 26056 5472
rect 25992 5412 25996 5468
rect 25996 5412 26052 5468
rect 26052 5412 26056 5468
rect 25992 5408 26056 5412
rect 3252 4924 3316 4928
rect 3252 4868 3256 4924
rect 3256 4868 3312 4924
rect 3312 4868 3316 4924
rect 3252 4864 3316 4868
rect 3332 4924 3396 4928
rect 3332 4868 3336 4924
rect 3336 4868 3392 4924
rect 3392 4868 3396 4924
rect 3332 4864 3396 4868
rect 3412 4924 3476 4928
rect 3412 4868 3416 4924
rect 3416 4868 3472 4924
rect 3472 4868 3476 4924
rect 3412 4864 3476 4868
rect 3492 4924 3556 4928
rect 3492 4868 3496 4924
rect 3496 4868 3552 4924
rect 3552 4868 3556 4924
rect 3492 4864 3556 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 6412 4924 6476 4928
rect 6412 4868 6416 4924
rect 6416 4868 6472 4924
rect 6472 4868 6476 4924
rect 6412 4864 6476 4868
rect 6492 4924 6556 4928
rect 6492 4868 6496 4924
rect 6496 4868 6552 4924
rect 6552 4868 6556 4924
rect 6492 4864 6556 4868
rect 9252 4924 9316 4928
rect 9252 4868 9256 4924
rect 9256 4868 9312 4924
rect 9312 4868 9316 4924
rect 9252 4864 9316 4868
rect 9332 4924 9396 4928
rect 9332 4868 9336 4924
rect 9336 4868 9392 4924
rect 9392 4868 9396 4924
rect 9332 4864 9396 4868
rect 9412 4924 9476 4928
rect 9412 4868 9416 4924
rect 9416 4868 9472 4924
rect 9472 4868 9476 4924
rect 9412 4864 9476 4868
rect 9492 4924 9556 4928
rect 9492 4868 9496 4924
rect 9496 4868 9552 4924
rect 9552 4868 9556 4924
rect 9492 4864 9556 4868
rect 12252 4924 12316 4928
rect 12252 4868 12256 4924
rect 12256 4868 12312 4924
rect 12312 4868 12316 4924
rect 12252 4864 12316 4868
rect 12332 4924 12396 4928
rect 12332 4868 12336 4924
rect 12336 4868 12392 4924
rect 12392 4868 12396 4924
rect 12332 4864 12396 4868
rect 12412 4924 12476 4928
rect 12412 4868 12416 4924
rect 12416 4868 12472 4924
rect 12472 4868 12476 4924
rect 12412 4864 12476 4868
rect 12492 4924 12556 4928
rect 12492 4868 12496 4924
rect 12496 4868 12552 4924
rect 12552 4868 12556 4924
rect 12492 4864 12556 4868
rect 15252 4924 15316 4928
rect 15252 4868 15256 4924
rect 15256 4868 15312 4924
rect 15312 4868 15316 4924
rect 15252 4864 15316 4868
rect 15332 4924 15396 4928
rect 15332 4868 15336 4924
rect 15336 4868 15392 4924
rect 15392 4868 15396 4924
rect 15332 4864 15396 4868
rect 15412 4924 15476 4928
rect 15412 4868 15416 4924
rect 15416 4868 15472 4924
rect 15472 4868 15476 4924
rect 15412 4864 15476 4868
rect 15492 4924 15556 4928
rect 15492 4868 15496 4924
rect 15496 4868 15552 4924
rect 15552 4868 15556 4924
rect 15492 4864 15556 4868
rect 18252 4924 18316 4928
rect 18252 4868 18256 4924
rect 18256 4868 18312 4924
rect 18312 4868 18316 4924
rect 18252 4864 18316 4868
rect 18332 4924 18396 4928
rect 18332 4868 18336 4924
rect 18336 4868 18392 4924
rect 18392 4868 18396 4924
rect 18332 4864 18396 4868
rect 18412 4924 18476 4928
rect 18412 4868 18416 4924
rect 18416 4868 18472 4924
rect 18472 4868 18476 4924
rect 18412 4864 18476 4868
rect 18492 4924 18556 4928
rect 18492 4868 18496 4924
rect 18496 4868 18552 4924
rect 18552 4868 18556 4924
rect 18492 4864 18556 4868
rect 21252 4924 21316 4928
rect 21252 4868 21256 4924
rect 21256 4868 21312 4924
rect 21312 4868 21316 4924
rect 21252 4864 21316 4868
rect 21332 4924 21396 4928
rect 21332 4868 21336 4924
rect 21336 4868 21392 4924
rect 21392 4868 21396 4924
rect 21332 4864 21396 4868
rect 21412 4924 21476 4928
rect 21412 4868 21416 4924
rect 21416 4868 21472 4924
rect 21472 4868 21476 4924
rect 21412 4864 21476 4868
rect 21492 4924 21556 4928
rect 21492 4868 21496 4924
rect 21496 4868 21552 4924
rect 21552 4868 21556 4924
rect 21492 4864 21556 4868
rect 24252 4924 24316 4928
rect 24252 4868 24256 4924
rect 24256 4868 24312 4924
rect 24312 4868 24316 4924
rect 24252 4864 24316 4868
rect 24332 4924 24396 4928
rect 24332 4868 24336 4924
rect 24336 4868 24392 4924
rect 24392 4868 24396 4924
rect 24332 4864 24396 4868
rect 24412 4924 24476 4928
rect 24412 4868 24416 4924
rect 24416 4868 24472 4924
rect 24472 4868 24476 4924
rect 24412 4864 24476 4868
rect 24492 4924 24556 4928
rect 24492 4868 24496 4924
rect 24496 4868 24552 4924
rect 24552 4868 24556 4924
rect 24492 4864 24556 4868
rect 27252 4924 27316 4928
rect 27252 4868 27256 4924
rect 27256 4868 27312 4924
rect 27312 4868 27316 4924
rect 27252 4864 27316 4868
rect 27332 4924 27396 4928
rect 27332 4868 27336 4924
rect 27336 4868 27392 4924
rect 27392 4868 27396 4924
rect 27332 4864 27396 4868
rect 27412 4924 27476 4928
rect 27412 4868 27416 4924
rect 27416 4868 27472 4924
rect 27472 4868 27476 4924
rect 27412 4864 27476 4868
rect 27492 4924 27556 4928
rect 27492 4868 27496 4924
rect 27496 4868 27552 4924
rect 27552 4868 27556 4924
rect 27492 4864 27556 4868
rect 1752 4380 1816 4384
rect 1752 4324 1756 4380
rect 1756 4324 1812 4380
rect 1812 4324 1816 4380
rect 1752 4320 1816 4324
rect 1832 4380 1896 4384
rect 1832 4324 1836 4380
rect 1836 4324 1892 4380
rect 1892 4324 1896 4380
rect 1832 4320 1896 4324
rect 1912 4380 1976 4384
rect 1912 4324 1916 4380
rect 1916 4324 1972 4380
rect 1972 4324 1976 4380
rect 1912 4320 1976 4324
rect 1992 4380 2056 4384
rect 1992 4324 1996 4380
rect 1996 4324 2052 4380
rect 2052 4324 2056 4380
rect 1992 4320 2056 4324
rect 4752 4380 4816 4384
rect 4752 4324 4756 4380
rect 4756 4324 4812 4380
rect 4812 4324 4816 4380
rect 4752 4320 4816 4324
rect 4832 4380 4896 4384
rect 4832 4324 4836 4380
rect 4836 4324 4892 4380
rect 4892 4324 4896 4380
rect 4832 4320 4896 4324
rect 4912 4380 4976 4384
rect 4912 4324 4916 4380
rect 4916 4324 4972 4380
rect 4972 4324 4976 4380
rect 4912 4320 4976 4324
rect 4992 4380 5056 4384
rect 4992 4324 4996 4380
rect 4996 4324 5052 4380
rect 5052 4324 5056 4380
rect 4992 4320 5056 4324
rect 7752 4380 7816 4384
rect 7752 4324 7756 4380
rect 7756 4324 7812 4380
rect 7812 4324 7816 4380
rect 7752 4320 7816 4324
rect 7832 4380 7896 4384
rect 7832 4324 7836 4380
rect 7836 4324 7892 4380
rect 7892 4324 7896 4380
rect 7832 4320 7896 4324
rect 7912 4380 7976 4384
rect 7912 4324 7916 4380
rect 7916 4324 7972 4380
rect 7972 4324 7976 4380
rect 7912 4320 7976 4324
rect 7992 4380 8056 4384
rect 7992 4324 7996 4380
rect 7996 4324 8052 4380
rect 8052 4324 8056 4380
rect 7992 4320 8056 4324
rect 10752 4380 10816 4384
rect 10752 4324 10756 4380
rect 10756 4324 10812 4380
rect 10812 4324 10816 4380
rect 10752 4320 10816 4324
rect 10832 4380 10896 4384
rect 10832 4324 10836 4380
rect 10836 4324 10892 4380
rect 10892 4324 10896 4380
rect 10832 4320 10896 4324
rect 10912 4380 10976 4384
rect 10912 4324 10916 4380
rect 10916 4324 10972 4380
rect 10972 4324 10976 4380
rect 10912 4320 10976 4324
rect 10992 4380 11056 4384
rect 10992 4324 10996 4380
rect 10996 4324 11052 4380
rect 11052 4324 11056 4380
rect 10992 4320 11056 4324
rect 13752 4380 13816 4384
rect 13752 4324 13756 4380
rect 13756 4324 13812 4380
rect 13812 4324 13816 4380
rect 13752 4320 13816 4324
rect 13832 4380 13896 4384
rect 13832 4324 13836 4380
rect 13836 4324 13892 4380
rect 13892 4324 13896 4380
rect 13832 4320 13896 4324
rect 13912 4380 13976 4384
rect 13912 4324 13916 4380
rect 13916 4324 13972 4380
rect 13972 4324 13976 4380
rect 13912 4320 13976 4324
rect 13992 4380 14056 4384
rect 13992 4324 13996 4380
rect 13996 4324 14052 4380
rect 14052 4324 14056 4380
rect 13992 4320 14056 4324
rect 16752 4380 16816 4384
rect 16752 4324 16756 4380
rect 16756 4324 16812 4380
rect 16812 4324 16816 4380
rect 16752 4320 16816 4324
rect 16832 4380 16896 4384
rect 16832 4324 16836 4380
rect 16836 4324 16892 4380
rect 16892 4324 16896 4380
rect 16832 4320 16896 4324
rect 16912 4380 16976 4384
rect 16912 4324 16916 4380
rect 16916 4324 16972 4380
rect 16972 4324 16976 4380
rect 16912 4320 16976 4324
rect 16992 4380 17056 4384
rect 16992 4324 16996 4380
rect 16996 4324 17052 4380
rect 17052 4324 17056 4380
rect 16992 4320 17056 4324
rect 19752 4380 19816 4384
rect 19752 4324 19756 4380
rect 19756 4324 19812 4380
rect 19812 4324 19816 4380
rect 19752 4320 19816 4324
rect 19832 4380 19896 4384
rect 19832 4324 19836 4380
rect 19836 4324 19892 4380
rect 19892 4324 19896 4380
rect 19832 4320 19896 4324
rect 19912 4380 19976 4384
rect 19912 4324 19916 4380
rect 19916 4324 19972 4380
rect 19972 4324 19976 4380
rect 19912 4320 19976 4324
rect 19992 4380 20056 4384
rect 19992 4324 19996 4380
rect 19996 4324 20052 4380
rect 20052 4324 20056 4380
rect 19992 4320 20056 4324
rect 22752 4380 22816 4384
rect 22752 4324 22756 4380
rect 22756 4324 22812 4380
rect 22812 4324 22816 4380
rect 22752 4320 22816 4324
rect 22832 4380 22896 4384
rect 22832 4324 22836 4380
rect 22836 4324 22892 4380
rect 22892 4324 22896 4380
rect 22832 4320 22896 4324
rect 22912 4380 22976 4384
rect 22912 4324 22916 4380
rect 22916 4324 22972 4380
rect 22972 4324 22976 4380
rect 22912 4320 22976 4324
rect 22992 4380 23056 4384
rect 22992 4324 22996 4380
rect 22996 4324 23052 4380
rect 23052 4324 23056 4380
rect 22992 4320 23056 4324
rect 25752 4380 25816 4384
rect 25752 4324 25756 4380
rect 25756 4324 25812 4380
rect 25812 4324 25816 4380
rect 25752 4320 25816 4324
rect 25832 4380 25896 4384
rect 25832 4324 25836 4380
rect 25836 4324 25892 4380
rect 25892 4324 25896 4380
rect 25832 4320 25896 4324
rect 25912 4380 25976 4384
rect 25912 4324 25916 4380
rect 25916 4324 25972 4380
rect 25972 4324 25976 4380
rect 25912 4320 25976 4324
rect 25992 4380 26056 4384
rect 25992 4324 25996 4380
rect 25996 4324 26052 4380
rect 26052 4324 26056 4380
rect 25992 4320 26056 4324
rect 3252 3836 3316 3840
rect 3252 3780 3256 3836
rect 3256 3780 3312 3836
rect 3312 3780 3316 3836
rect 3252 3776 3316 3780
rect 3332 3836 3396 3840
rect 3332 3780 3336 3836
rect 3336 3780 3392 3836
rect 3392 3780 3396 3836
rect 3332 3776 3396 3780
rect 3412 3836 3476 3840
rect 3412 3780 3416 3836
rect 3416 3780 3472 3836
rect 3472 3780 3476 3836
rect 3412 3776 3476 3780
rect 3492 3836 3556 3840
rect 3492 3780 3496 3836
rect 3496 3780 3552 3836
rect 3552 3780 3556 3836
rect 3492 3776 3556 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 6412 3836 6476 3840
rect 6412 3780 6416 3836
rect 6416 3780 6472 3836
rect 6472 3780 6476 3836
rect 6412 3776 6476 3780
rect 6492 3836 6556 3840
rect 6492 3780 6496 3836
rect 6496 3780 6552 3836
rect 6552 3780 6556 3836
rect 6492 3776 6556 3780
rect 9252 3836 9316 3840
rect 9252 3780 9256 3836
rect 9256 3780 9312 3836
rect 9312 3780 9316 3836
rect 9252 3776 9316 3780
rect 9332 3836 9396 3840
rect 9332 3780 9336 3836
rect 9336 3780 9392 3836
rect 9392 3780 9396 3836
rect 9332 3776 9396 3780
rect 9412 3836 9476 3840
rect 9412 3780 9416 3836
rect 9416 3780 9472 3836
rect 9472 3780 9476 3836
rect 9412 3776 9476 3780
rect 9492 3836 9556 3840
rect 9492 3780 9496 3836
rect 9496 3780 9552 3836
rect 9552 3780 9556 3836
rect 9492 3776 9556 3780
rect 12252 3836 12316 3840
rect 12252 3780 12256 3836
rect 12256 3780 12312 3836
rect 12312 3780 12316 3836
rect 12252 3776 12316 3780
rect 12332 3836 12396 3840
rect 12332 3780 12336 3836
rect 12336 3780 12392 3836
rect 12392 3780 12396 3836
rect 12332 3776 12396 3780
rect 12412 3836 12476 3840
rect 12412 3780 12416 3836
rect 12416 3780 12472 3836
rect 12472 3780 12476 3836
rect 12412 3776 12476 3780
rect 12492 3836 12556 3840
rect 12492 3780 12496 3836
rect 12496 3780 12552 3836
rect 12552 3780 12556 3836
rect 12492 3776 12556 3780
rect 15252 3836 15316 3840
rect 15252 3780 15256 3836
rect 15256 3780 15312 3836
rect 15312 3780 15316 3836
rect 15252 3776 15316 3780
rect 15332 3836 15396 3840
rect 15332 3780 15336 3836
rect 15336 3780 15392 3836
rect 15392 3780 15396 3836
rect 15332 3776 15396 3780
rect 15412 3836 15476 3840
rect 15412 3780 15416 3836
rect 15416 3780 15472 3836
rect 15472 3780 15476 3836
rect 15412 3776 15476 3780
rect 15492 3836 15556 3840
rect 15492 3780 15496 3836
rect 15496 3780 15552 3836
rect 15552 3780 15556 3836
rect 15492 3776 15556 3780
rect 18252 3836 18316 3840
rect 18252 3780 18256 3836
rect 18256 3780 18312 3836
rect 18312 3780 18316 3836
rect 18252 3776 18316 3780
rect 18332 3836 18396 3840
rect 18332 3780 18336 3836
rect 18336 3780 18392 3836
rect 18392 3780 18396 3836
rect 18332 3776 18396 3780
rect 18412 3836 18476 3840
rect 18412 3780 18416 3836
rect 18416 3780 18472 3836
rect 18472 3780 18476 3836
rect 18412 3776 18476 3780
rect 18492 3836 18556 3840
rect 18492 3780 18496 3836
rect 18496 3780 18552 3836
rect 18552 3780 18556 3836
rect 18492 3776 18556 3780
rect 21252 3836 21316 3840
rect 21252 3780 21256 3836
rect 21256 3780 21312 3836
rect 21312 3780 21316 3836
rect 21252 3776 21316 3780
rect 21332 3836 21396 3840
rect 21332 3780 21336 3836
rect 21336 3780 21392 3836
rect 21392 3780 21396 3836
rect 21332 3776 21396 3780
rect 21412 3836 21476 3840
rect 21412 3780 21416 3836
rect 21416 3780 21472 3836
rect 21472 3780 21476 3836
rect 21412 3776 21476 3780
rect 21492 3836 21556 3840
rect 21492 3780 21496 3836
rect 21496 3780 21552 3836
rect 21552 3780 21556 3836
rect 21492 3776 21556 3780
rect 24252 3836 24316 3840
rect 24252 3780 24256 3836
rect 24256 3780 24312 3836
rect 24312 3780 24316 3836
rect 24252 3776 24316 3780
rect 24332 3836 24396 3840
rect 24332 3780 24336 3836
rect 24336 3780 24392 3836
rect 24392 3780 24396 3836
rect 24332 3776 24396 3780
rect 24412 3836 24476 3840
rect 24412 3780 24416 3836
rect 24416 3780 24472 3836
rect 24472 3780 24476 3836
rect 24412 3776 24476 3780
rect 24492 3836 24556 3840
rect 24492 3780 24496 3836
rect 24496 3780 24552 3836
rect 24552 3780 24556 3836
rect 24492 3776 24556 3780
rect 27252 3836 27316 3840
rect 27252 3780 27256 3836
rect 27256 3780 27312 3836
rect 27312 3780 27316 3836
rect 27252 3776 27316 3780
rect 27332 3836 27396 3840
rect 27332 3780 27336 3836
rect 27336 3780 27392 3836
rect 27392 3780 27396 3836
rect 27332 3776 27396 3780
rect 27412 3836 27476 3840
rect 27412 3780 27416 3836
rect 27416 3780 27472 3836
rect 27472 3780 27476 3836
rect 27412 3776 27476 3780
rect 27492 3836 27556 3840
rect 27492 3780 27496 3836
rect 27496 3780 27552 3836
rect 27552 3780 27556 3836
rect 27492 3776 27556 3780
rect 1752 3292 1816 3296
rect 1752 3236 1756 3292
rect 1756 3236 1812 3292
rect 1812 3236 1816 3292
rect 1752 3232 1816 3236
rect 1832 3292 1896 3296
rect 1832 3236 1836 3292
rect 1836 3236 1892 3292
rect 1892 3236 1896 3292
rect 1832 3232 1896 3236
rect 1912 3292 1976 3296
rect 1912 3236 1916 3292
rect 1916 3236 1972 3292
rect 1972 3236 1976 3292
rect 1912 3232 1976 3236
rect 1992 3292 2056 3296
rect 1992 3236 1996 3292
rect 1996 3236 2052 3292
rect 2052 3236 2056 3292
rect 1992 3232 2056 3236
rect 4752 3292 4816 3296
rect 4752 3236 4756 3292
rect 4756 3236 4812 3292
rect 4812 3236 4816 3292
rect 4752 3232 4816 3236
rect 4832 3292 4896 3296
rect 4832 3236 4836 3292
rect 4836 3236 4892 3292
rect 4892 3236 4896 3292
rect 4832 3232 4896 3236
rect 4912 3292 4976 3296
rect 4912 3236 4916 3292
rect 4916 3236 4972 3292
rect 4972 3236 4976 3292
rect 4912 3232 4976 3236
rect 4992 3292 5056 3296
rect 4992 3236 4996 3292
rect 4996 3236 5052 3292
rect 5052 3236 5056 3292
rect 4992 3232 5056 3236
rect 7752 3292 7816 3296
rect 7752 3236 7756 3292
rect 7756 3236 7812 3292
rect 7812 3236 7816 3292
rect 7752 3232 7816 3236
rect 7832 3292 7896 3296
rect 7832 3236 7836 3292
rect 7836 3236 7892 3292
rect 7892 3236 7896 3292
rect 7832 3232 7896 3236
rect 7912 3292 7976 3296
rect 7912 3236 7916 3292
rect 7916 3236 7972 3292
rect 7972 3236 7976 3292
rect 7912 3232 7976 3236
rect 7992 3292 8056 3296
rect 7992 3236 7996 3292
rect 7996 3236 8052 3292
rect 8052 3236 8056 3292
rect 7992 3232 8056 3236
rect 10752 3292 10816 3296
rect 10752 3236 10756 3292
rect 10756 3236 10812 3292
rect 10812 3236 10816 3292
rect 10752 3232 10816 3236
rect 10832 3292 10896 3296
rect 10832 3236 10836 3292
rect 10836 3236 10892 3292
rect 10892 3236 10896 3292
rect 10832 3232 10896 3236
rect 10912 3292 10976 3296
rect 10912 3236 10916 3292
rect 10916 3236 10972 3292
rect 10972 3236 10976 3292
rect 10912 3232 10976 3236
rect 10992 3292 11056 3296
rect 10992 3236 10996 3292
rect 10996 3236 11052 3292
rect 11052 3236 11056 3292
rect 10992 3232 11056 3236
rect 13752 3292 13816 3296
rect 13752 3236 13756 3292
rect 13756 3236 13812 3292
rect 13812 3236 13816 3292
rect 13752 3232 13816 3236
rect 13832 3292 13896 3296
rect 13832 3236 13836 3292
rect 13836 3236 13892 3292
rect 13892 3236 13896 3292
rect 13832 3232 13896 3236
rect 13912 3292 13976 3296
rect 13912 3236 13916 3292
rect 13916 3236 13972 3292
rect 13972 3236 13976 3292
rect 13912 3232 13976 3236
rect 13992 3292 14056 3296
rect 13992 3236 13996 3292
rect 13996 3236 14052 3292
rect 14052 3236 14056 3292
rect 13992 3232 14056 3236
rect 16752 3292 16816 3296
rect 16752 3236 16756 3292
rect 16756 3236 16812 3292
rect 16812 3236 16816 3292
rect 16752 3232 16816 3236
rect 16832 3292 16896 3296
rect 16832 3236 16836 3292
rect 16836 3236 16892 3292
rect 16892 3236 16896 3292
rect 16832 3232 16896 3236
rect 16912 3292 16976 3296
rect 16912 3236 16916 3292
rect 16916 3236 16972 3292
rect 16972 3236 16976 3292
rect 16912 3232 16976 3236
rect 16992 3292 17056 3296
rect 16992 3236 16996 3292
rect 16996 3236 17052 3292
rect 17052 3236 17056 3292
rect 16992 3232 17056 3236
rect 19752 3292 19816 3296
rect 19752 3236 19756 3292
rect 19756 3236 19812 3292
rect 19812 3236 19816 3292
rect 19752 3232 19816 3236
rect 19832 3292 19896 3296
rect 19832 3236 19836 3292
rect 19836 3236 19892 3292
rect 19892 3236 19896 3292
rect 19832 3232 19896 3236
rect 19912 3292 19976 3296
rect 19912 3236 19916 3292
rect 19916 3236 19972 3292
rect 19972 3236 19976 3292
rect 19912 3232 19976 3236
rect 19992 3292 20056 3296
rect 19992 3236 19996 3292
rect 19996 3236 20052 3292
rect 20052 3236 20056 3292
rect 19992 3232 20056 3236
rect 22752 3292 22816 3296
rect 22752 3236 22756 3292
rect 22756 3236 22812 3292
rect 22812 3236 22816 3292
rect 22752 3232 22816 3236
rect 22832 3292 22896 3296
rect 22832 3236 22836 3292
rect 22836 3236 22892 3292
rect 22892 3236 22896 3292
rect 22832 3232 22896 3236
rect 22912 3292 22976 3296
rect 22912 3236 22916 3292
rect 22916 3236 22972 3292
rect 22972 3236 22976 3292
rect 22912 3232 22976 3236
rect 22992 3292 23056 3296
rect 22992 3236 22996 3292
rect 22996 3236 23052 3292
rect 23052 3236 23056 3292
rect 22992 3232 23056 3236
rect 25752 3292 25816 3296
rect 25752 3236 25756 3292
rect 25756 3236 25812 3292
rect 25812 3236 25816 3292
rect 25752 3232 25816 3236
rect 25832 3292 25896 3296
rect 25832 3236 25836 3292
rect 25836 3236 25892 3292
rect 25892 3236 25896 3292
rect 25832 3232 25896 3236
rect 25912 3292 25976 3296
rect 25912 3236 25916 3292
rect 25916 3236 25972 3292
rect 25972 3236 25976 3292
rect 25912 3232 25976 3236
rect 25992 3292 26056 3296
rect 25992 3236 25996 3292
rect 25996 3236 26052 3292
rect 26052 3236 26056 3292
rect 25992 3232 26056 3236
rect 3252 2748 3316 2752
rect 3252 2692 3256 2748
rect 3256 2692 3312 2748
rect 3312 2692 3316 2748
rect 3252 2688 3316 2692
rect 3332 2748 3396 2752
rect 3332 2692 3336 2748
rect 3336 2692 3392 2748
rect 3392 2692 3396 2748
rect 3332 2688 3396 2692
rect 3412 2748 3476 2752
rect 3412 2692 3416 2748
rect 3416 2692 3472 2748
rect 3472 2692 3476 2748
rect 3412 2688 3476 2692
rect 3492 2748 3556 2752
rect 3492 2692 3496 2748
rect 3496 2692 3552 2748
rect 3552 2692 3556 2748
rect 3492 2688 3556 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 6412 2748 6476 2752
rect 6412 2692 6416 2748
rect 6416 2692 6472 2748
rect 6472 2692 6476 2748
rect 6412 2688 6476 2692
rect 6492 2748 6556 2752
rect 6492 2692 6496 2748
rect 6496 2692 6552 2748
rect 6552 2692 6556 2748
rect 6492 2688 6556 2692
rect 9252 2748 9316 2752
rect 9252 2692 9256 2748
rect 9256 2692 9312 2748
rect 9312 2692 9316 2748
rect 9252 2688 9316 2692
rect 9332 2748 9396 2752
rect 9332 2692 9336 2748
rect 9336 2692 9392 2748
rect 9392 2692 9396 2748
rect 9332 2688 9396 2692
rect 9412 2748 9476 2752
rect 9412 2692 9416 2748
rect 9416 2692 9472 2748
rect 9472 2692 9476 2748
rect 9412 2688 9476 2692
rect 9492 2748 9556 2752
rect 9492 2692 9496 2748
rect 9496 2692 9552 2748
rect 9552 2692 9556 2748
rect 9492 2688 9556 2692
rect 12252 2748 12316 2752
rect 12252 2692 12256 2748
rect 12256 2692 12312 2748
rect 12312 2692 12316 2748
rect 12252 2688 12316 2692
rect 12332 2748 12396 2752
rect 12332 2692 12336 2748
rect 12336 2692 12392 2748
rect 12392 2692 12396 2748
rect 12332 2688 12396 2692
rect 12412 2748 12476 2752
rect 12412 2692 12416 2748
rect 12416 2692 12472 2748
rect 12472 2692 12476 2748
rect 12412 2688 12476 2692
rect 12492 2748 12556 2752
rect 12492 2692 12496 2748
rect 12496 2692 12552 2748
rect 12552 2692 12556 2748
rect 12492 2688 12556 2692
rect 15252 2748 15316 2752
rect 15252 2692 15256 2748
rect 15256 2692 15312 2748
rect 15312 2692 15316 2748
rect 15252 2688 15316 2692
rect 15332 2748 15396 2752
rect 15332 2692 15336 2748
rect 15336 2692 15392 2748
rect 15392 2692 15396 2748
rect 15332 2688 15396 2692
rect 15412 2748 15476 2752
rect 15412 2692 15416 2748
rect 15416 2692 15472 2748
rect 15472 2692 15476 2748
rect 15412 2688 15476 2692
rect 15492 2748 15556 2752
rect 15492 2692 15496 2748
rect 15496 2692 15552 2748
rect 15552 2692 15556 2748
rect 15492 2688 15556 2692
rect 18252 2748 18316 2752
rect 18252 2692 18256 2748
rect 18256 2692 18312 2748
rect 18312 2692 18316 2748
rect 18252 2688 18316 2692
rect 18332 2748 18396 2752
rect 18332 2692 18336 2748
rect 18336 2692 18392 2748
rect 18392 2692 18396 2748
rect 18332 2688 18396 2692
rect 18412 2748 18476 2752
rect 18412 2692 18416 2748
rect 18416 2692 18472 2748
rect 18472 2692 18476 2748
rect 18412 2688 18476 2692
rect 18492 2748 18556 2752
rect 18492 2692 18496 2748
rect 18496 2692 18552 2748
rect 18552 2692 18556 2748
rect 18492 2688 18556 2692
rect 21252 2748 21316 2752
rect 21252 2692 21256 2748
rect 21256 2692 21312 2748
rect 21312 2692 21316 2748
rect 21252 2688 21316 2692
rect 21332 2748 21396 2752
rect 21332 2692 21336 2748
rect 21336 2692 21392 2748
rect 21392 2692 21396 2748
rect 21332 2688 21396 2692
rect 21412 2748 21476 2752
rect 21412 2692 21416 2748
rect 21416 2692 21472 2748
rect 21472 2692 21476 2748
rect 21412 2688 21476 2692
rect 21492 2748 21556 2752
rect 21492 2692 21496 2748
rect 21496 2692 21552 2748
rect 21552 2692 21556 2748
rect 21492 2688 21556 2692
rect 24252 2748 24316 2752
rect 24252 2692 24256 2748
rect 24256 2692 24312 2748
rect 24312 2692 24316 2748
rect 24252 2688 24316 2692
rect 24332 2748 24396 2752
rect 24332 2692 24336 2748
rect 24336 2692 24392 2748
rect 24392 2692 24396 2748
rect 24332 2688 24396 2692
rect 24412 2748 24476 2752
rect 24412 2692 24416 2748
rect 24416 2692 24472 2748
rect 24472 2692 24476 2748
rect 24412 2688 24476 2692
rect 24492 2748 24556 2752
rect 24492 2692 24496 2748
rect 24496 2692 24552 2748
rect 24552 2692 24556 2748
rect 24492 2688 24556 2692
rect 27252 2748 27316 2752
rect 27252 2692 27256 2748
rect 27256 2692 27312 2748
rect 27312 2692 27316 2748
rect 27252 2688 27316 2692
rect 27332 2748 27396 2752
rect 27332 2692 27336 2748
rect 27336 2692 27392 2748
rect 27392 2692 27396 2748
rect 27332 2688 27396 2692
rect 27412 2748 27476 2752
rect 27412 2692 27416 2748
rect 27416 2692 27472 2748
rect 27472 2692 27476 2748
rect 27412 2688 27476 2692
rect 27492 2748 27556 2752
rect 27492 2692 27496 2748
rect 27496 2692 27552 2748
rect 27552 2692 27556 2748
rect 27492 2688 27556 2692
rect 1752 2204 1816 2208
rect 1752 2148 1756 2204
rect 1756 2148 1812 2204
rect 1812 2148 1816 2204
rect 1752 2144 1816 2148
rect 1832 2204 1896 2208
rect 1832 2148 1836 2204
rect 1836 2148 1892 2204
rect 1892 2148 1896 2204
rect 1832 2144 1896 2148
rect 1912 2204 1976 2208
rect 1912 2148 1916 2204
rect 1916 2148 1972 2204
rect 1972 2148 1976 2204
rect 1912 2144 1976 2148
rect 1992 2204 2056 2208
rect 1992 2148 1996 2204
rect 1996 2148 2052 2204
rect 2052 2148 2056 2204
rect 1992 2144 2056 2148
rect 4752 2204 4816 2208
rect 4752 2148 4756 2204
rect 4756 2148 4812 2204
rect 4812 2148 4816 2204
rect 4752 2144 4816 2148
rect 4832 2204 4896 2208
rect 4832 2148 4836 2204
rect 4836 2148 4892 2204
rect 4892 2148 4896 2204
rect 4832 2144 4896 2148
rect 4912 2204 4976 2208
rect 4912 2148 4916 2204
rect 4916 2148 4972 2204
rect 4972 2148 4976 2204
rect 4912 2144 4976 2148
rect 4992 2204 5056 2208
rect 4992 2148 4996 2204
rect 4996 2148 5052 2204
rect 5052 2148 5056 2204
rect 4992 2144 5056 2148
rect 7752 2204 7816 2208
rect 7752 2148 7756 2204
rect 7756 2148 7812 2204
rect 7812 2148 7816 2204
rect 7752 2144 7816 2148
rect 7832 2204 7896 2208
rect 7832 2148 7836 2204
rect 7836 2148 7892 2204
rect 7892 2148 7896 2204
rect 7832 2144 7896 2148
rect 7912 2204 7976 2208
rect 7912 2148 7916 2204
rect 7916 2148 7972 2204
rect 7972 2148 7976 2204
rect 7912 2144 7976 2148
rect 7992 2204 8056 2208
rect 7992 2148 7996 2204
rect 7996 2148 8052 2204
rect 8052 2148 8056 2204
rect 7992 2144 8056 2148
rect 10752 2204 10816 2208
rect 10752 2148 10756 2204
rect 10756 2148 10812 2204
rect 10812 2148 10816 2204
rect 10752 2144 10816 2148
rect 10832 2204 10896 2208
rect 10832 2148 10836 2204
rect 10836 2148 10892 2204
rect 10892 2148 10896 2204
rect 10832 2144 10896 2148
rect 10912 2204 10976 2208
rect 10912 2148 10916 2204
rect 10916 2148 10972 2204
rect 10972 2148 10976 2204
rect 10912 2144 10976 2148
rect 10992 2204 11056 2208
rect 10992 2148 10996 2204
rect 10996 2148 11052 2204
rect 11052 2148 11056 2204
rect 10992 2144 11056 2148
rect 13752 2204 13816 2208
rect 13752 2148 13756 2204
rect 13756 2148 13812 2204
rect 13812 2148 13816 2204
rect 13752 2144 13816 2148
rect 13832 2204 13896 2208
rect 13832 2148 13836 2204
rect 13836 2148 13892 2204
rect 13892 2148 13896 2204
rect 13832 2144 13896 2148
rect 13912 2204 13976 2208
rect 13912 2148 13916 2204
rect 13916 2148 13972 2204
rect 13972 2148 13976 2204
rect 13912 2144 13976 2148
rect 13992 2204 14056 2208
rect 13992 2148 13996 2204
rect 13996 2148 14052 2204
rect 14052 2148 14056 2204
rect 13992 2144 14056 2148
rect 16752 2204 16816 2208
rect 16752 2148 16756 2204
rect 16756 2148 16812 2204
rect 16812 2148 16816 2204
rect 16752 2144 16816 2148
rect 16832 2204 16896 2208
rect 16832 2148 16836 2204
rect 16836 2148 16892 2204
rect 16892 2148 16896 2204
rect 16832 2144 16896 2148
rect 16912 2204 16976 2208
rect 16912 2148 16916 2204
rect 16916 2148 16972 2204
rect 16972 2148 16976 2204
rect 16912 2144 16976 2148
rect 16992 2204 17056 2208
rect 16992 2148 16996 2204
rect 16996 2148 17052 2204
rect 17052 2148 17056 2204
rect 16992 2144 17056 2148
rect 19752 2204 19816 2208
rect 19752 2148 19756 2204
rect 19756 2148 19812 2204
rect 19812 2148 19816 2204
rect 19752 2144 19816 2148
rect 19832 2204 19896 2208
rect 19832 2148 19836 2204
rect 19836 2148 19892 2204
rect 19892 2148 19896 2204
rect 19832 2144 19896 2148
rect 19912 2204 19976 2208
rect 19912 2148 19916 2204
rect 19916 2148 19972 2204
rect 19972 2148 19976 2204
rect 19912 2144 19976 2148
rect 19992 2204 20056 2208
rect 19992 2148 19996 2204
rect 19996 2148 20052 2204
rect 20052 2148 20056 2204
rect 19992 2144 20056 2148
rect 22752 2204 22816 2208
rect 22752 2148 22756 2204
rect 22756 2148 22812 2204
rect 22812 2148 22816 2204
rect 22752 2144 22816 2148
rect 22832 2204 22896 2208
rect 22832 2148 22836 2204
rect 22836 2148 22892 2204
rect 22892 2148 22896 2204
rect 22832 2144 22896 2148
rect 22912 2204 22976 2208
rect 22912 2148 22916 2204
rect 22916 2148 22972 2204
rect 22972 2148 22976 2204
rect 22912 2144 22976 2148
rect 22992 2204 23056 2208
rect 22992 2148 22996 2204
rect 22996 2148 23052 2204
rect 23052 2148 23056 2204
rect 22992 2144 23056 2148
rect 25752 2204 25816 2208
rect 25752 2148 25756 2204
rect 25756 2148 25812 2204
rect 25812 2148 25816 2204
rect 25752 2144 25816 2148
rect 25832 2204 25896 2208
rect 25832 2148 25836 2204
rect 25836 2148 25892 2204
rect 25892 2148 25896 2204
rect 25832 2144 25896 2148
rect 25912 2204 25976 2208
rect 25912 2148 25916 2204
rect 25916 2148 25972 2204
rect 25972 2148 25976 2204
rect 25912 2144 25976 2148
rect 25992 2204 26056 2208
rect 25992 2148 25996 2204
rect 25996 2148 26052 2204
rect 26052 2148 26056 2204
rect 25992 2144 26056 2148
<< metal4 >>
rect 1744 29408 2064 29424
rect 1744 29344 1752 29408
rect 1816 29344 1832 29408
rect 1896 29344 1912 29408
rect 1976 29344 1992 29408
rect 2056 29344 2064 29408
rect 1744 28320 2064 29344
rect 1744 28256 1752 28320
rect 1816 28256 1832 28320
rect 1896 28256 1912 28320
rect 1976 28256 1992 28320
rect 2056 28256 2064 28320
rect 1744 27232 2064 28256
rect 1744 27168 1752 27232
rect 1816 27168 1832 27232
rect 1896 27168 1912 27232
rect 1976 27168 1992 27232
rect 2056 27168 2064 27232
rect 1744 27046 2064 27168
rect 1744 26810 1786 27046
rect 2022 26810 2064 27046
rect 1744 26144 2064 26810
rect 1744 26080 1752 26144
rect 1816 26080 1832 26144
rect 1896 26080 1912 26144
rect 1976 26080 1992 26144
rect 2056 26080 2064 26144
rect 1744 25056 2064 26080
rect 1744 24992 1752 25056
rect 1816 24992 1832 25056
rect 1896 24992 1912 25056
rect 1976 24992 1992 25056
rect 2056 24992 2064 25056
rect 1744 24046 2064 24992
rect 1744 23968 1786 24046
rect 2022 23968 2064 24046
rect 1744 23904 1752 23968
rect 2056 23904 2064 23968
rect 1744 23810 1786 23904
rect 2022 23810 2064 23904
rect 1744 22880 2064 23810
rect 1744 22816 1752 22880
rect 1816 22816 1832 22880
rect 1896 22816 1912 22880
rect 1976 22816 1992 22880
rect 2056 22816 2064 22880
rect 1744 21792 2064 22816
rect 1744 21728 1752 21792
rect 1816 21728 1832 21792
rect 1896 21728 1912 21792
rect 1976 21728 1992 21792
rect 2056 21728 2064 21792
rect 1744 21046 2064 21728
rect 1744 20810 1786 21046
rect 2022 20810 2064 21046
rect 1744 20704 2064 20810
rect 1744 20640 1752 20704
rect 1816 20640 1832 20704
rect 1896 20640 1912 20704
rect 1976 20640 1992 20704
rect 2056 20640 2064 20704
rect 1744 19616 2064 20640
rect 1744 19552 1752 19616
rect 1816 19552 1832 19616
rect 1896 19552 1912 19616
rect 1976 19552 1992 19616
rect 2056 19552 2064 19616
rect 1744 18528 2064 19552
rect 1744 18464 1752 18528
rect 1816 18464 1832 18528
rect 1896 18464 1912 18528
rect 1976 18464 1992 18528
rect 2056 18464 2064 18528
rect 1744 18046 2064 18464
rect 1744 17810 1786 18046
rect 2022 17810 2064 18046
rect 1744 17440 2064 17810
rect 1744 17376 1752 17440
rect 1816 17376 1832 17440
rect 1896 17376 1912 17440
rect 1976 17376 1992 17440
rect 2056 17376 2064 17440
rect 1744 16352 2064 17376
rect 1744 16288 1752 16352
rect 1816 16288 1832 16352
rect 1896 16288 1912 16352
rect 1976 16288 1992 16352
rect 2056 16288 2064 16352
rect 1744 15264 2064 16288
rect 1744 15200 1752 15264
rect 1816 15200 1832 15264
rect 1896 15200 1912 15264
rect 1976 15200 1992 15264
rect 2056 15200 2064 15264
rect 1744 15046 2064 15200
rect 1744 14810 1786 15046
rect 2022 14810 2064 15046
rect 1744 14176 2064 14810
rect 1744 14112 1752 14176
rect 1816 14112 1832 14176
rect 1896 14112 1912 14176
rect 1976 14112 1992 14176
rect 2056 14112 2064 14176
rect 1744 13088 2064 14112
rect 1744 13024 1752 13088
rect 1816 13024 1832 13088
rect 1896 13024 1912 13088
rect 1976 13024 1992 13088
rect 2056 13024 2064 13088
rect 1744 12046 2064 13024
rect 1744 12000 1786 12046
rect 2022 12000 2064 12046
rect 1744 11936 1752 12000
rect 2056 11936 2064 12000
rect 1744 11810 1786 11936
rect 2022 11810 2064 11936
rect 1744 10912 2064 11810
rect 1744 10848 1752 10912
rect 1816 10848 1832 10912
rect 1896 10848 1912 10912
rect 1976 10848 1992 10912
rect 2056 10848 2064 10912
rect 1744 9824 2064 10848
rect 1744 9760 1752 9824
rect 1816 9760 1832 9824
rect 1896 9760 1912 9824
rect 1976 9760 1992 9824
rect 2056 9760 2064 9824
rect 1744 9046 2064 9760
rect 1744 8810 1786 9046
rect 2022 8810 2064 9046
rect 1744 8736 2064 8810
rect 1744 8672 1752 8736
rect 1816 8672 1832 8736
rect 1896 8672 1912 8736
rect 1976 8672 1992 8736
rect 2056 8672 2064 8736
rect 1744 7648 2064 8672
rect 1744 7584 1752 7648
rect 1816 7584 1832 7648
rect 1896 7584 1912 7648
rect 1976 7584 1992 7648
rect 2056 7584 2064 7648
rect 1744 6560 2064 7584
rect 1744 6496 1752 6560
rect 1816 6496 1832 6560
rect 1896 6496 1912 6560
rect 1976 6496 1992 6560
rect 2056 6496 2064 6560
rect 1744 6046 2064 6496
rect 1744 5810 1786 6046
rect 2022 5810 2064 6046
rect 1744 5472 2064 5810
rect 1744 5408 1752 5472
rect 1816 5408 1832 5472
rect 1896 5408 1912 5472
rect 1976 5408 1992 5472
rect 2056 5408 2064 5472
rect 1744 4384 2064 5408
rect 1744 4320 1752 4384
rect 1816 4320 1832 4384
rect 1896 4320 1912 4384
rect 1976 4320 1992 4384
rect 2056 4320 2064 4384
rect 1744 3296 2064 4320
rect 1744 3232 1752 3296
rect 1816 3232 1832 3296
rect 1896 3232 1912 3296
rect 1976 3232 1992 3296
rect 2056 3232 2064 3296
rect 1744 3046 2064 3232
rect 1744 2810 1786 3046
rect 2022 2810 2064 3046
rect 1744 2208 2064 2810
rect 1744 2144 1752 2208
rect 1816 2144 1832 2208
rect 1896 2144 1912 2208
rect 1976 2144 1992 2208
rect 2056 2144 2064 2208
rect 1744 2128 2064 2144
rect 3244 28864 3564 29424
rect 3244 28800 3252 28864
rect 3316 28800 3332 28864
rect 3396 28800 3412 28864
rect 3476 28800 3492 28864
rect 3556 28800 3564 28864
rect 3244 28546 3564 28800
rect 3244 28310 3286 28546
rect 3522 28310 3564 28546
rect 3244 27776 3564 28310
rect 3244 27712 3252 27776
rect 3316 27712 3332 27776
rect 3396 27712 3412 27776
rect 3476 27712 3492 27776
rect 3556 27712 3564 27776
rect 3244 26688 3564 27712
rect 3244 26624 3252 26688
rect 3316 26624 3332 26688
rect 3396 26624 3412 26688
rect 3476 26624 3492 26688
rect 3556 26624 3564 26688
rect 3244 25600 3564 26624
rect 3244 25536 3252 25600
rect 3316 25546 3332 25600
rect 3396 25546 3412 25600
rect 3476 25546 3492 25600
rect 3556 25536 3564 25600
rect 3244 25310 3286 25536
rect 3522 25310 3564 25536
rect 3244 24512 3564 25310
rect 3244 24448 3252 24512
rect 3316 24448 3332 24512
rect 3396 24448 3412 24512
rect 3476 24448 3492 24512
rect 3556 24448 3564 24512
rect 3244 23424 3564 24448
rect 3244 23360 3252 23424
rect 3316 23360 3332 23424
rect 3396 23360 3412 23424
rect 3476 23360 3492 23424
rect 3556 23360 3564 23424
rect 3244 22546 3564 23360
rect 3244 22336 3286 22546
rect 3522 22336 3564 22546
rect 3244 22272 3252 22336
rect 3316 22272 3332 22310
rect 3396 22272 3412 22310
rect 3476 22272 3492 22310
rect 3556 22272 3564 22336
rect 3244 21248 3564 22272
rect 3244 21184 3252 21248
rect 3316 21184 3332 21248
rect 3396 21184 3412 21248
rect 3476 21184 3492 21248
rect 3556 21184 3564 21248
rect 3244 20160 3564 21184
rect 3244 20096 3252 20160
rect 3316 20096 3332 20160
rect 3396 20096 3412 20160
rect 3476 20096 3492 20160
rect 3556 20096 3564 20160
rect 3244 19546 3564 20096
rect 3244 19310 3286 19546
rect 3522 19310 3564 19546
rect 3244 19072 3564 19310
rect 3244 19008 3252 19072
rect 3316 19008 3332 19072
rect 3396 19008 3412 19072
rect 3476 19008 3492 19072
rect 3556 19008 3564 19072
rect 3244 17984 3564 19008
rect 3244 17920 3252 17984
rect 3316 17920 3332 17984
rect 3396 17920 3412 17984
rect 3476 17920 3492 17984
rect 3556 17920 3564 17984
rect 3244 16896 3564 17920
rect 3244 16832 3252 16896
rect 3316 16832 3332 16896
rect 3396 16832 3412 16896
rect 3476 16832 3492 16896
rect 3556 16832 3564 16896
rect 3244 16546 3564 16832
rect 3244 16310 3286 16546
rect 3522 16310 3564 16546
rect 3244 15808 3564 16310
rect 3244 15744 3252 15808
rect 3316 15744 3332 15808
rect 3396 15744 3412 15808
rect 3476 15744 3492 15808
rect 3556 15744 3564 15808
rect 3244 14720 3564 15744
rect 3244 14656 3252 14720
rect 3316 14656 3332 14720
rect 3396 14656 3412 14720
rect 3476 14656 3492 14720
rect 3556 14656 3564 14720
rect 3244 13632 3564 14656
rect 3244 13568 3252 13632
rect 3316 13568 3332 13632
rect 3396 13568 3412 13632
rect 3476 13568 3492 13632
rect 3556 13568 3564 13632
rect 3244 13546 3564 13568
rect 3244 13310 3286 13546
rect 3522 13310 3564 13546
rect 3244 12544 3564 13310
rect 3244 12480 3252 12544
rect 3316 12480 3332 12544
rect 3396 12480 3412 12544
rect 3476 12480 3492 12544
rect 3556 12480 3564 12544
rect 3244 11456 3564 12480
rect 3244 11392 3252 11456
rect 3316 11392 3332 11456
rect 3396 11392 3412 11456
rect 3476 11392 3492 11456
rect 3556 11392 3564 11456
rect 3244 10546 3564 11392
rect 3244 10368 3286 10546
rect 3522 10368 3564 10546
rect 3244 10304 3252 10368
rect 3316 10304 3332 10310
rect 3396 10304 3412 10310
rect 3476 10304 3492 10310
rect 3556 10304 3564 10368
rect 3244 9280 3564 10304
rect 3244 9216 3252 9280
rect 3316 9216 3332 9280
rect 3396 9216 3412 9280
rect 3476 9216 3492 9280
rect 3556 9216 3564 9280
rect 3244 8192 3564 9216
rect 3244 8128 3252 8192
rect 3316 8128 3332 8192
rect 3396 8128 3412 8192
rect 3476 8128 3492 8192
rect 3556 8128 3564 8192
rect 3244 7546 3564 8128
rect 3244 7310 3286 7546
rect 3522 7310 3564 7546
rect 3244 7104 3564 7310
rect 3244 7040 3252 7104
rect 3316 7040 3332 7104
rect 3396 7040 3412 7104
rect 3476 7040 3492 7104
rect 3556 7040 3564 7104
rect 3244 6016 3564 7040
rect 3244 5952 3252 6016
rect 3316 5952 3332 6016
rect 3396 5952 3412 6016
rect 3476 5952 3492 6016
rect 3556 5952 3564 6016
rect 3244 4928 3564 5952
rect 3244 4864 3252 4928
rect 3316 4864 3332 4928
rect 3396 4864 3412 4928
rect 3476 4864 3492 4928
rect 3556 4864 3564 4928
rect 3244 4546 3564 4864
rect 3244 4310 3286 4546
rect 3522 4310 3564 4546
rect 3244 3840 3564 4310
rect 3244 3776 3252 3840
rect 3316 3776 3332 3840
rect 3396 3776 3412 3840
rect 3476 3776 3492 3840
rect 3556 3776 3564 3840
rect 3244 2752 3564 3776
rect 3244 2688 3252 2752
rect 3316 2688 3332 2752
rect 3396 2688 3412 2752
rect 3476 2688 3492 2752
rect 3556 2688 3564 2752
rect 3244 2128 3564 2688
rect 4744 29408 5064 29424
rect 4744 29344 4752 29408
rect 4816 29344 4832 29408
rect 4896 29344 4912 29408
rect 4976 29344 4992 29408
rect 5056 29344 5064 29408
rect 4744 28320 5064 29344
rect 4744 28256 4752 28320
rect 4816 28256 4832 28320
rect 4896 28256 4912 28320
rect 4976 28256 4992 28320
rect 5056 28256 5064 28320
rect 4744 27232 5064 28256
rect 4744 27168 4752 27232
rect 4816 27168 4832 27232
rect 4896 27168 4912 27232
rect 4976 27168 4992 27232
rect 5056 27168 5064 27232
rect 4744 27046 5064 27168
rect 4744 26810 4786 27046
rect 5022 26810 5064 27046
rect 4744 26144 5064 26810
rect 4744 26080 4752 26144
rect 4816 26080 4832 26144
rect 4896 26080 4912 26144
rect 4976 26080 4992 26144
rect 5056 26080 5064 26144
rect 4744 25056 5064 26080
rect 4744 24992 4752 25056
rect 4816 24992 4832 25056
rect 4896 24992 4912 25056
rect 4976 24992 4992 25056
rect 5056 24992 5064 25056
rect 4744 24046 5064 24992
rect 4744 23968 4786 24046
rect 5022 23968 5064 24046
rect 4744 23904 4752 23968
rect 5056 23904 5064 23968
rect 4744 23810 4786 23904
rect 5022 23810 5064 23904
rect 4744 22880 5064 23810
rect 4744 22816 4752 22880
rect 4816 22816 4832 22880
rect 4896 22816 4912 22880
rect 4976 22816 4992 22880
rect 5056 22816 5064 22880
rect 4744 21792 5064 22816
rect 4744 21728 4752 21792
rect 4816 21728 4832 21792
rect 4896 21728 4912 21792
rect 4976 21728 4992 21792
rect 5056 21728 5064 21792
rect 4744 21046 5064 21728
rect 4744 20810 4786 21046
rect 5022 20810 5064 21046
rect 4744 20704 5064 20810
rect 4744 20640 4752 20704
rect 4816 20640 4832 20704
rect 4896 20640 4912 20704
rect 4976 20640 4992 20704
rect 5056 20640 5064 20704
rect 4744 19616 5064 20640
rect 4744 19552 4752 19616
rect 4816 19552 4832 19616
rect 4896 19552 4912 19616
rect 4976 19552 4992 19616
rect 5056 19552 5064 19616
rect 4744 18528 5064 19552
rect 4744 18464 4752 18528
rect 4816 18464 4832 18528
rect 4896 18464 4912 18528
rect 4976 18464 4992 18528
rect 5056 18464 5064 18528
rect 4744 18046 5064 18464
rect 4744 17810 4786 18046
rect 5022 17810 5064 18046
rect 4744 17440 5064 17810
rect 4744 17376 4752 17440
rect 4816 17376 4832 17440
rect 4896 17376 4912 17440
rect 4976 17376 4992 17440
rect 5056 17376 5064 17440
rect 4744 16352 5064 17376
rect 4744 16288 4752 16352
rect 4816 16288 4832 16352
rect 4896 16288 4912 16352
rect 4976 16288 4992 16352
rect 5056 16288 5064 16352
rect 4744 15264 5064 16288
rect 4744 15200 4752 15264
rect 4816 15200 4832 15264
rect 4896 15200 4912 15264
rect 4976 15200 4992 15264
rect 5056 15200 5064 15264
rect 4744 15046 5064 15200
rect 4744 14810 4786 15046
rect 5022 14810 5064 15046
rect 4744 14176 5064 14810
rect 4744 14112 4752 14176
rect 4816 14112 4832 14176
rect 4896 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5064 14176
rect 4744 13088 5064 14112
rect 4744 13024 4752 13088
rect 4816 13024 4832 13088
rect 4896 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5064 13088
rect 4744 12046 5064 13024
rect 4744 12000 4786 12046
rect 5022 12000 5064 12046
rect 4744 11936 4752 12000
rect 5056 11936 5064 12000
rect 4744 11810 4786 11936
rect 5022 11810 5064 11936
rect 4744 10912 5064 11810
rect 4744 10848 4752 10912
rect 4816 10848 4832 10912
rect 4896 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5064 10912
rect 4744 9824 5064 10848
rect 4744 9760 4752 9824
rect 4816 9760 4832 9824
rect 4896 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5064 9824
rect 4744 9046 5064 9760
rect 4744 8810 4786 9046
rect 5022 8810 5064 9046
rect 4744 8736 5064 8810
rect 4744 8672 4752 8736
rect 4816 8672 4832 8736
rect 4896 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5064 8736
rect 4744 7648 5064 8672
rect 4744 7584 4752 7648
rect 4816 7584 4832 7648
rect 4896 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5064 7648
rect 4744 6560 5064 7584
rect 4744 6496 4752 6560
rect 4816 6496 4832 6560
rect 4896 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5064 6560
rect 4744 6046 5064 6496
rect 4744 5810 4786 6046
rect 5022 5810 5064 6046
rect 4744 5472 5064 5810
rect 4744 5408 4752 5472
rect 4816 5408 4832 5472
rect 4896 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5064 5472
rect 4744 4384 5064 5408
rect 4744 4320 4752 4384
rect 4816 4320 4832 4384
rect 4896 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5064 4384
rect 4744 3296 5064 4320
rect 4744 3232 4752 3296
rect 4816 3232 4832 3296
rect 4896 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5064 3296
rect 4744 3046 5064 3232
rect 4744 2810 4786 3046
rect 5022 2810 5064 3046
rect 4744 2208 5064 2810
rect 4744 2144 4752 2208
rect 4816 2144 4832 2208
rect 4896 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5064 2208
rect 4744 2128 5064 2144
rect 6244 28864 6564 29424
rect 6244 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6412 28864
rect 6476 28800 6492 28864
rect 6556 28800 6564 28864
rect 6244 28546 6564 28800
rect 6244 28310 6286 28546
rect 6522 28310 6564 28546
rect 6244 27776 6564 28310
rect 6244 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6412 27776
rect 6476 27712 6492 27776
rect 6556 27712 6564 27776
rect 6244 26688 6564 27712
rect 6244 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6412 26688
rect 6476 26624 6492 26688
rect 6556 26624 6564 26688
rect 6244 25600 6564 26624
rect 6244 25536 6252 25600
rect 6316 25546 6332 25600
rect 6396 25546 6412 25600
rect 6476 25546 6492 25600
rect 6556 25536 6564 25600
rect 6244 25310 6286 25536
rect 6522 25310 6564 25536
rect 6244 24512 6564 25310
rect 6244 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6412 24512
rect 6476 24448 6492 24512
rect 6556 24448 6564 24512
rect 6244 23424 6564 24448
rect 6244 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6412 23424
rect 6476 23360 6492 23424
rect 6556 23360 6564 23424
rect 6244 22546 6564 23360
rect 6244 22336 6286 22546
rect 6522 22336 6564 22546
rect 6244 22272 6252 22336
rect 6316 22272 6332 22310
rect 6396 22272 6412 22310
rect 6476 22272 6492 22310
rect 6556 22272 6564 22336
rect 6244 21248 6564 22272
rect 6244 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6412 21248
rect 6476 21184 6492 21248
rect 6556 21184 6564 21248
rect 6244 20160 6564 21184
rect 6244 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6412 20160
rect 6476 20096 6492 20160
rect 6556 20096 6564 20160
rect 6244 19546 6564 20096
rect 6244 19310 6286 19546
rect 6522 19310 6564 19546
rect 6244 19072 6564 19310
rect 6244 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6412 19072
rect 6476 19008 6492 19072
rect 6556 19008 6564 19072
rect 6244 17984 6564 19008
rect 6244 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6412 17984
rect 6476 17920 6492 17984
rect 6556 17920 6564 17984
rect 6244 16896 6564 17920
rect 6244 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6412 16896
rect 6476 16832 6492 16896
rect 6556 16832 6564 16896
rect 6244 16546 6564 16832
rect 6244 16310 6286 16546
rect 6522 16310 6564 16546
rect 6244 15808 6564 16310
rect 6244 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6412 15808
rect 6476 15744 6492 15808
rect 6556 15744 6564 15808
rect 6244 14720 6564 15744
rect 6244 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6412 14720
rect 6476 14656 6492 14720
rect 6556 14656 6564 14720
rect 6244 13632 6564 14656
rect 6244 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6412 13632
rect 6476 13568 6492 13632
rect 6556 13568 6564 13632
rect 6244 13546 6564 13568
rect 6244 13310 6286 13546
rect 6522 13310 6564 13546
rect 6244 12544 6564 13310
rect 6244 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6412 12544
rect 6476 12480 6492 12544
rect 6556 12480 6564 12544
rect 6244 11456 6564 12480
rect 6244 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6412 11456
rect 6476 11392 6492 11456
rect 6556 11392 6564 11456
rect 6244 10546 6564 11392
rect 6244 10368 6286 10546
rect 6522 10368 6564 10546
rect 6244 10304 6252 10368
rect 6316 10304 6332 10310
rect 6396 10304 6412 10310
rect 6476 10304 6492 10310
rect 6556 10304 6564 10368
rect 6244 9280 6564 10304
rect 6244 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6412 9280
rect 6476 9216 6492 9280
rect 6556 9216 6564 9280
rect 6244 8192 6564 9216
rect 6244 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6412 8192
rect 6476 8128 6492 8192
rect 6556 8128 6564 8192
rect 6244 7546 6564 8128
rect 6244 7310 6286 7546
rect 6522 7310 6564 7546
rect 6244 7104 6564 7310
rect 6244 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6412 7104
rect 6476 7040 6492 7104
rect 6556 7040 6564 7104
rect 6244 6016 6564 7040
rect 6244 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6412 6016
rect 6476 5952 6492 6016
rect 6556 5952 6564 6016
rect 6244 4928 6564 5952
rect 6244 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6412 4928
rect 6476 4864 6492 4928
rect 6556 4864 6564 4928
rect 6244 4546 6564 4864
rect 6244 4310 6286 4546
rect 6522 4310 6564 4546
rect 6244 3840 6564 4310
rect 6244 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6412 3840
rect 6476 3776 6492 3840
rect 6556 3776 6564 3840
rect 6244 2752 6564 3776
rect 6244 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6412 2752
rect 6476 2688 6492 2752
rect 6556 2688 6564 2752
rect 6244 2128 6564 2688
rect 7744 29408 8064 29424
rect 7744 29344 7752 29408
rect 7816 29344 7832 29408
rect 7896 29344 7912 29408
rect 7976 29344 7992 29408
rect 8056 29344 8064 29408
rect 7744 28320 8064 29344
rect 7744 28256 7752 28320
rect 7816 28256 7832 28320
rect 7896 28256 7912 28320
rect 7976 28256 7992 28320
rect 8056 28256 8064 28320
rect 7744 27232 8064 28256
rect 7744 27168 7752 27232
rect 7816 27168 7832 27232
rect 7896 27168 7912 27232
rect 7976 27168 7992 27232
rect 8056 27168 8064 27232
rect 7744 27046 8064 27168
rect 7744 26810 7786 27046
rect 8022 26810 8064 27046
rect 7744 26144 8064 26810
rect 7744 26080 7752 26144
rect 7816 26080 7832 26144
rect 7896 26080 7912 26144
rect 7976 26080 7992 26144
rect 8056 26080 8064 26144
rect 7744 25056 8064 26080
rect 7744 24992 7752 25056
rect 7816 24992 7832 25056
rect 7896 24992 7912 25056
rect 7976 24992 7992 25056
rect 8056 24992 8064 25056
rect 7744 24046 8064 24992
rect 7744 23968 7786 24046
rect 8022 23968 8064 24046
rect 7744 23904 7752 23968
rect 8056 23904 8064 23968
rect 7744 23810 7786 23904
rect 8022 23810 8064 23904
rect 7744 22880 8064 23810
rect 7744 22816 7752 22880
rect 7816 22816 7832 22880
rect 7896 22816 7912 22880
rect 7976 22816 7992 22880
rect 8056 22816 8064 22880
rect 7744 21792 8064 22816
rect 7744 21728 7752 21792
rect 7816 21728 7832 21792
rect 7896 21728 7912 21792
rect 7976 21728 7992 21792
rect 8056 21728 8064 21792
rect 7744 21046 8064 21728
rect 7744 20810 7786 21046
rect 8022 20810 8064 21046
rect 7744 20704 8064 20810
rect 7744 20640 7752 20704
rect 7816 20640 7832 20704
rect 7896 20640 7912 20704
rect 7976 20640 7992 20704
rect 8056 20640 8064 20704
rect 7744 19616 8064 20640
rect 7744 19552 7752 19616
rect 7816 19552 7832 19616
rect 7896 19552 7912 19616
rect 7976 19552 7992 19616
rect 8056 19552 8064 19616
rect 7744 18528 8064 19552
rect 7744 18464 7752 18528
rect 7816 18464 7832 18528
rect 7896 18464 7912 18528
rect 7976 18464 7992 18528
rect 8056 18464 8064 18528
rect 7744 18046 8064 18464
rect 7744 17810 7786 18046
rect 8022 17810 8064 18046
rect 7744 17440 8064 17810
rect 7744 17376 7752 17440
rect 7816 17376 7832 17440
rect 7896 17376 7912 17440
rect 7976 17376 7992 17440
rect 8056 17376 8064 17440
rect 7744 16352 8064 17376
rect 7744 16288 7752 16352
rect 7816 16288 7832 16352
rect 7896 16288 7912 16352
rect 7976 16288 7992 16352
rect 8056 16288 8064 16352
rect 7744 15264 8064 16288
rect 7744 15200 7752 15264
rect 7816 15200 7832 15264
rect 7896 15200 7912 15264
rect 7976 15200 7992 15264
rect 8056 15200 8064 15264
rect 7744 15046 8064 15200
rect 7744 14810 7786 15046
rect 8022 14810 8064 15046
rect 7744 14176 8064 14810
rect 7744 14112 7752 14176
rect 7816 14112 7832 14176
rect 7896 14112 7912 14176
rect 7976 14112 7992 14176
rect 8056 14112 8064 14176
rect 7744 13088 8064 14112
rect 7744 13024 7752 13088
rect 7816 13024 7832 13088
rect 7896 13024 7912 13088
rect 7976 13024 7992 13088
rect 8056 13024 8064 13088
rect 7744 12046 8064 13024
rect 7744 12000 7786 12046
rect 8022 12000 8064 12046
rect 7744 11936 7752 12000
rect 8056 11936 8064 12000
rect 7744 11810 7786 11936
rect 8022 11810 8064 11936
rect 7744 10912 8064 11810
rect 7744 10848 7752 10912
rect 7816 10848 7832 10912
rect 7896 10848 7912 10912
rect 7976 10848 7992 10912
rect 8056 10848 8064 10912
rect 7744 9824 8064 10848
rect 7744 9760 7752 9824
rect 7816 9760 7832 9824
rect 7896 9760 7912 9824
rect 7976 9760 7992 9824
rect 8056 9760 8064 9824
rect 7744 9046 8064 9760
rect 7744 8810 7786 9046
rect 8022 8810 8064 9046
rect 7744 8736 8064 8810
rect 7744 8672 7752 8736
rect 7816 8672 7832 8736
rect 7896 8672 7912 8736
rect 7976 8672 7992 8736
rect 8056 8672 8064 8736
rect 7744 7648 8064 8672
rect 7744 7584 7752 7648
rect 7816 7584 7832 7648
rect 7896 7584 7912 7648
rect 7976 7584 7992 7648
rect 8056 7584 8064 7648
rect 7744 6560 8064 7584
rect 7744 6496 7752 6560
rect 7816 6496 7832 6560
rect 7896 6496 7912 6560
rect 7976 6496 7992 6560
rect 8056 6496 8064 6560
rect 7744 6046 8064 6496
rect 7744 5810 7786 6046
rect 8022 5810 8064 6046
rect 7744 5472 8064 5810
rect 7744 5408 7752 5472
rect 7816 5408 7832 5472
rect 7896 5408 7912 5472
rect 7976 5408 7992 5472
rect 8056 5408 8064 5472
rect 7744 4384 8064 5408
rect 7744 4320 7752 4384
rect 7816 4320 7832 4384
rect 7896 4320 7912 4384
rect 7976 4320 7992 4384
rect 8056 4320 8064 4384
rect 7744 3296 8064 4320
rect 7744 3232 7752 3296
rect 7816 3232 7832 3296
rect 7896 3232 7912 3296
rect 7976 3232 7992 3296
rect 8056 3232 8064 3296
rect 7744 3046 8064 3232
rect 7744 2810 7786 3046
rect 8022 2810 8064 3046
rect 7744 2208 8064 2810
rect 7744 2144 7752 2208
rect 7816 2144 7832 2208
rect 7896 2144 7912 2208
rect 7976 2144 7992 2208
rect 8056 2144 8064 2208
rect 7744 2128 8064 2144
rect 9244 28864 9564 29424
rect 9244 28800 9252 28864
rect 9316 28800 9332 28864
rect 9396 28800 9412 28864
rect 9476 28800 9492 28864
rect 9556 28800 9564 28864
rect 9244 28546 9564 28800
rect 9244 28310 9286 28546
rect 9522 28310 9564 28546
rect 9244 27776 9564 28310
rect 9244 27712 9252 27776
rect 9316 27712 9332 27776
rect 9396 27712 9412 27776
rect 9476 27712 9492 27776
rect 9556 27712 9564 27776
rect 9244 26688 9564 27712
rect 9244 26624 9252 26688
rect 9316 26624 9332 26688
rect 9396 26624 9412 26688
rect 9476 26624 9492 26688
rect 9556 26624 9564 26688
rect 9244 25600 9564 26624
rect 9244 25536 9252 25600
rect 9316 25546 9332 25600
rect 9396 25546 9412 25600
rect 9476 25546 9492 25600
rect 9556 25536 9564 25600
rect 9244 25310 9286 25536
rect 9522 25310 9564 25536
rect 9244 24512 9564 25310
rect 9244 24448 9252 24512
rect 9316 24448 9332 24512
rect 9396 24448 9412 24512
rect 9476 24448 9492 24512
rect 9556 24448 9564 24512
rect 9244 23424 9564 24448
rect 9244 23360 9252 23424
rect 9316 23360 9332 23424
rect 9396 23360 9412 23424
rect 9476 23360 9492 23424
rect 9556 23360 9564 23424
rect 9244 22546 9564 23360
rect 9244 22336 9286 22546
rect 9522 22336 9564 22546
rect 9244 22272 9252 22336
rect 9316 22272 9332 22310
rect 9396 22272 9412 22310
rect 9476 22272 9492 22310
rect 9556 22272 9564 22336
rect 9244 21248 9564 22272
rect 9244 21184 9252 21248
rect 9316 21184 9332 21248
rect 9396 21184 9412 21248
rect 9476 21184 9492 21248
rect 9556 21184 9564 21248
rect 9244 20160 9564 21184
rect 9244 20096 9252 20160
rect 9316 20096 9332 20160
rect 9396 20096 9412 20160
rect 9476 20096 9492 20160
rect 9556 20096 9564 20160
rect 9244 19546 9564 20096
rect 9244 19310 9286 19546
rect 9522 19310 9564 19546
rect 9244 19072 9564 19310
rect 9244 19008 9252 19072
rect 9316 19008 9332 19072
rect 9396 19008 9412 19072
rect 9476 19008 9492 19072
rect 9556 19008 9564 19072
rect 9244 17984 9564 19008
rect 9244 17920 9252 17984
rect 9316 17920 9332 17984
rect 9396 17920 9412 17984
rect 9476 17920 9492 17984
rect 9556 17920 9564 17984
rect 9244 16896 9564 17920
rect 9244 16832 9252 16896
rect 9316 16832 9332 16896
rect 9396 16832 9412 16896
rect 9476 16832 9492 16896
rect 9556 16832 9564 16896
rect 9244 16546 9564 16832
rect 9244 16310 9286 16546
rect 9522 16310 9564 16546
rect 9244 15808 9564 16310
rect 9244 15744 9252 15808
rect 9316 15744 9332 15808
rect 9396 15744 9412 15808
rect 9476 15744 9492 15808
rect 9556 15744 9564 15808
rect 9244 14720 9564 15744
rect 9244 14656 9252 14720
rect 9316 14656 9332 14720
rect 9396 14656 9412 14720
rect 9476 14656 9492 14720
rect 9556 14656 9564 14720
rect 9244 13632 9564 14656
rect 9244 13568 9252 13632
rect 9316 13568 9332 13632
rect 9396 13568 9412 13632
rect 9476 13568 9492 13632
rect 9556 13568 9564 13632
rect 9244 13546 9564 13568
rect 9244 13310 9286 13546
rect 9522 13310 9564 13546
rect 9244 12544 9564 13310
rect 9244 12480 9252 12544
rect 9316 12480 9332 12544
rect 9396 12480 9412 12544
rect 9476 12480 9492 12544
rect 9556 12480 9564 12544
rect 9244 11456 9564 12480
rect 9244 11392 9252 11456
rect 9316 11392 9332 11456
rect 9396 11392 9412 11456
rect 9476 11392 9492 11456
rect 9556 11392 9564 11456
rect 9244 10546 9564 11392
rect 9244 10368 9286 10546
rect 9522 10368 9564 10546
rect 9244 10304 9252 10368
rect 9316 10304 9332 10310
rect 9396 10304 9412 10310
rect 9476 10304 9492 10310
rect 9556 10304 9564 10368
rect 9244 9280 9564 10304
rect 9244 9216 9252 9280
rect 9316 9216 9332 9280
rect 9396 9216 9412 9280
rect 9476 9216 9492 9280
rect 9556 9216 9564 9280
rect 9244 8192 9564 9216
rect 9244 8128 9252 8192
rect 9316 8128 9332 8192
rect 9396 8128 9412 8192
rect 9476 8128 9492 8192
rect 9556 8128 9564 8192
rect 9244 7546 9564 8128
rect 9244 7310 9286 7546
rect 9522 7310 9564 7546
rect 9244 7104 9564 7310
rect 9244 7040 9252 7104
rect 9316 7040 9332 7104
rect 9396 7040 9412 7104
rect 9476 7040 9492 7104
rect 9556 7040 9564 7104
rect 9244 6016 9564 7040
rect 9244 5952 9252 6016
rect 9316 5952 9332 6016
rect 9396 5952 9412 6016
rect 9476 5952 9492 6016
rect 9556 5952 9564 6016
rect 9244 4928 9564 5952
rect 9244 4864 9252 4928
rect 9316 4864 9332 4928
rect 9396 4864 9412 4928
rect 9476 4864 9492 4928
rect 9556 4864 9564 4928
rect 9244 4546 9564 4864
rect 9244 4310 9286 4546
rect 9522 4310 9564 4546
rect 9244 3840 9564 4310
rect 9244 3776 9252 3840
rect 9316 3776 9332 3840
rect 9396 3776 9412 3840
rect 9476 3776 9492 3840
rect 9556 3776 9564 3840
rect 9244 2752 9564 3776
rect 9244 2688 9252 2752
rect 9316 2688 9332 2752
rect 9396 2688 9412 2752
rect 9476 2688 9492 2752
rect 9556 2688 9564 2752
rect 9244 2128 9564 2688
rect 10744 29408 11064 29424
rect 10744 29344 10752 29408
rect 10816 29344 10832 29408
rect 10896 29344 10912 29408
rect 10976 29344 10992 29408
rect 11056 29344 11064 29408
rect 10744 28320 11064 29344
rect 10744 28256 10752 28320
rect 10816 28256 10832 28320
rect 10896 28256 10912 28320
rect 10976 28256 10992 28320
rect 11056 28256 11064 28320
rect 10744 27232 11064 28256
rect 10744 27168 10752 27232
rect 10816 27168 10832 27232
rect 10896 27168 10912 27232
rect 10976 27168 10992 27232
rect 11056 27168 11064 27232
rect 10744 27046 11064 27168
rect 10744 26810 10786 27046
rect 11022 26810 11064 27046
rect 10744 26144 11064 26810
rect 10744 26080 10752 26144
rect 10816 26080 10832 26144
rect 10896 26080 10912 26144
rect 10976 26080 10992 26144
rect 11056 26080 11064 26144
rect 10744 25056 11064 26080
rect 10744 24992 10752 25056
rect 10816 24992 10832 25056
rect 10896 24992 10912 25056
rect 10976 24992 10992 25056
rect 11056 24992 11064 25056
rect 10744 24046 11064 24992
rect 10744 23968 10786 24046
rect 11022 23968 11064 24046
rect 10744 23904 10752 23968
rect 11056 23904 11064 23968
rect 10744 23810 10786 23904
rect 11022 23810 11064 23904
rect 10744 22880 11064 23810
rect 10744 22816 10752 22880
rect 10816 22816 10832 22880
rect 10896 22816 10912 22880
rect 10976 22816 10992 22880
rect 11056 22816 11064 22880
rect 10744 21792 11064 22816
rect 10744 21728 10752 21792
rect 10816 21728 10832 21792
rect 10896 21728 10912 21792
rect 10976 21728 10992 21792
rect 11056 21728 11064 21792
rect 10744 21046 11064 21728
rect 10744 20810 10786 21046
rect 11022 20810 11064 21046
rect 10744 20704 11064 20810
rect 10744 20640 10752 20704
rect 10816 20640 10832 20704
rect 10896 20640 10912 20704
rect 10976 20640 10992 20704
rect 11056 20640 11064 20704
rect 10744 19616 11064 20640
rect 10744 19552 10752 19616
rect 10816 19552 10832 19616
rect 10896 19552 10912 19616
rect 10976 19552 10992 19616
rect 11056 19552 11064 19616
rect 10744 18528 11064 19552
rect 10744 18464 10752 18528
rect 10816 18464 10832 18528
rect 10896 18464 10912 18528
rect 10976 18464 10992 18528
rect 11056 18464 11064 18528
rect 10744 18046 11064 18464
rect 10744 17810 10786 18046
rect 11022 17810 11064 18046
rect 10744 17440 11064 17810
rect 10744 17376 10752 17440
rect 10816 17376 10832 17440
rect 10896 17376 10912 17440
rect 10976 17376 10992 17440
rect 11056 17376 11064 17440
rect 10744 16352 11064 17376
rect 10744 16288 10752 16352
rect 10816 16288 10832 16352
rect 10896 16288 10912 16352
rect 10976 16288 10992 16352
rect 11056 16288 11064 16352
rect 10744 15264 11064 16288
rect 10744 15200 10752 15264
rect 10816 15200 10832 15264
rect 10896 15200 10912 15264
rect 10976 15200 10992 15264
rect 11056 15200 11064 15264
rect 10744 15046 11064 15200
rect 10744 14810 10786 15046
rect 11022 14810 11064 15046
rect 10744 14176 11064 14810
rect 10744 14112 10752 14176
rect 10816 14112 10832 14176
rect 10896 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11064 14176
rect 10744 13088 11064 14112
rect 10744 13024 10752 13088
rect 10816 13024 10832 13088
rect 10896 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11064 13088
rect 10744 12046 11064 13024
rect 10744 12000 10786 12046
rect 11022 12000 11064 12046
rect 10744 11936 10752 12000
rect 11056 11936 11064 12000
rect 10744 11810 10786 11936
rect 11022 11810 11064 11936
rect 10744 10912 11064 11810
rect 10744 10848 10752 10912
rect 10816 10848 10832 10912
rect 10896 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11064 10912
rect 10744 9824 11064 10848
rect 10744 9760 10752 9824
rect 10816 9760 10832 9824
rect 10896 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11064 9824
rect 10744 9046 11064 9760
rect 10744 8810 10786 9046
rect 11022 8810 11064 9046
rect 10744 8736 11064 8810
rect 10744 8672 10752 8736
rect 10816 8672 10832 8736
rect 10896 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11064 8736
rect 10744 7648 11064 8672
rect 10744 7584 10752 7648
rect 10816 7584 10832 7648
rect 10896 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11064 7648
rect 10744 6560 11064 7584
rect 10744 6496 10752 6560
rect 10816 6496 10832 6560
rect 10896 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11064 6560
rect 10744 6046 11064 6496
rect 10744 5810 10786 6046
rect 11022 5810 11064 6046
rect 10744 5472 11064 5810
rect 10744 5408 10752 5472
rect 10816 5408 10832 5472
rect 10896 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11064 5472
rect 10744 4384 11064 5408
rect 10744 4320 10752 4384
rect 10816 4320 10832 4384
rect 10896 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11064 4384
rect 10744 3296 11064 4320
rect 10744 3232 10752 3296
rect 10816 3232 10832 3296
rect 10896 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11064 3296
rect 10744 3046 11064 3232
rect 10744 2810 10786 3046
rect 11022 2810 11064 3046
rect 10744 2208 11064 2810
rect 10744 2144 10752 2208
rect 10816 2144 10832 2208
rect 10896 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11064 2208
rect 10744 2128 11064 2144
rect 12244 28864 12564 29424
rect 12244 28800 12252 28864
rect 12316 28800 12332 28864
rect 12396 28800 12412 28864
rect 12476 28800 12492 28864
rect 12556 28800 12564 28864
rect 12244 28546 12564 28800
rect 12244 28310 12286 28546
rect 12522 28310 12564 28546
rect 12244 27776 12564 28310
rect 12244 27712 12252 27776
rect 12316 27712 12332 27776
rect 12396 27712 12412 27776
rect 12476 27712 12492 27776
rect 12556 27712 12564 27776
rect 12244 26688 12564 27712
rect 12244 26624 12252 26688
rect 12316 26624 12332 26688
rect 12396 26624 12412 26688
rect 12476 26624 12492 26688
rect 12556 26624 12564 26688
rect 12244 25600 12564 26624
rect 12244 25536 12252 25600
rect 12316 25546 12332 25600
rect 12396 25546 12412 25600
rect 12476 25546 12492 25600
rect 12556 25536 12564 25600
rect 12244 25310 12286 25536
rect 12522 25310 12564 25536
rect 12244 24512 12564 25310
rect 12244 24448 12252 24512
rect 12316 24448 12332 24512
rect 12396 24448 12412 24512
rect 12476 24448 12492 24512
rect 12556 24448 12564 24512
rect 12244 23424 12564 24448
rect 12244 23360 12252 23424
rect 12316 23360 12332 23424
rect 12396 23360 12412 23424
rect 12476 23360 12492 23424
rect 12556 23360 12564 23424
rect 12244 22546 12564 23360
rect 12244 22336 12286 22546
rect 12522 22336 12564 22546
rect 12244 22272 12252 22336
rect 12316 22272 12332 22310
rect 12396 22272 12412 22310
rect 12476 22272 12492 22310
rect 12556 22272 12564 22336
rect 12244 21248 12564 22272
rect 12244 21184 12252 21248
rect 12316 21184 12332 21248
rect 12396 21184 12412 21248
rect 12476 21184 12492 21248
rect 12556 21184 12564 21248
rect 12244 20160 12564 21184
rect 12244 20096 12252 20160
rect 12316 20096 12332 20160
rect 12396 20096 12412 20160
rect 12476 20096 12492 20160
rect 12556 20096 12564 20160
rect 12244 19546 12564 20096
rect 12244 19310 12286 19546
rect 12522 19310 12564 19546
rect 12244 19072 12564 19310
rect 12244 19008 12252 19072
rect 12316 19008 12332 19072
rect 12396 19008 12412 19072
rect 12476 19008 12492 19072
rect 12556 19008 12564 19072
rect 12244 17984 12564 19008
rect 12244 17920 12252 17984
rect 12316 17920 12332 17984
rect 12396 17920 12412 17984
rect 12476 17920 12492 17984
rect 12556 17920 12564 17984
rect 12244 16896 12564 17920
rect 12244 16832 12252 16896
rect 12316 16832 12332 16896
rect 12396 16832 12412 16896
rect 12476 16832 12492 16896
rect 12556 16832 12564 16896
rect 12244 16546 12564 16832
rect 12244 16310 12286 16546
rect 12522 16310 12564 16546
rect 12244 15808 12564 16310
rect 12244 15744 12252 15808
rect 12316 15744 12332 15808
rect 12396 15744 12412 15808
rect 12476 15744 12492 15808
rect 12556 15744 12564 15808
rect 12244 14720 12564 15744
rect 12244 14656 12252 14720
rect 12316 14656 12332 14720
rect 12396 14656 12412 14720
rect 12476 14656 12492 14720
rect 12556 14656 12564 14720
rect 12244 13632 12564 14656
rect 12244 13568 12252 13632
rect 12316 13568 12332 13632
rect 12396 13568 12412 13632
rect 12476 13568 12492 13632
rect 12556 13568 12564 13632
rect 12244 13546 12564 13568
rect 12244 13310 12286 13546
rect 12522 13310 12564 13546
rect 12244 12544 12564 13310
rect 12244 12480 12252 12544
rect 12316 12480 12332 12544
rect 12396 12480 12412 12544
rect 12476 12480 12492 12544
rect 12556 12480 12564 12544
rect 12244 11456 12564 12480
rect 12244 11392 12252 11456
rect 12316 11392 12332 11456
rect 12396 11392 12412 11456
rect 12476 11392 12492 11456
rect 12556 11392 12564 11456
rect 12244 10546 12564 11392
rect 12244 10368 12286 10546
rect 12522 10368 12564 10546
rect 12244 10304 12252 10368
rect 12316 10304 12332 10310
rect 12396 10304 12412 10310
rect 12476 10304 12492 10310
rect 12556 10304 12564 10368
rect 12244 9280 12564 10304
rect 12244 9216 12252 9280
rect 12316 9216 12332 9280
rect 12396 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12564 9280
rect 12244 8192 12564 9216
rect 12244 8128 12252 8192
rect 12316 8128 12332 8192
rect 12396 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12564 8192
rect 12244 7546 12564 8128
rect 12244 7310 12286 7546
rect 12522 7310 12564 7546
rect 12244 7104 12564 7310
rect 12244 7040 12252 7104
rect 12316 7040 12332 7104
rect 12396 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12564 7104
rect 12244 6016 12564 7040
rect 12244 5952 12252 6016
rect 12316 5952 12332 6016
rect 12396 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12564 6016
rect 12244 4928 12564 5952
rect 12244 4864 12252 4928
rect 12316 4864 12332 4928
rect 12396 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12564 4928
rect 12244 4546 12564 4864
rect 12244 4310 12286 4546
rect 12522 4310 12564 4546
rect 12244 3840 12564 4310
rect 12244 3776 12252 3840
rect 12316 3776 12332 3840
rect 12396 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12564 3840
rect 12244 2752 12564 3776
rect 12244 2688 12252 2752
rect 12316 2688 12332 2752
rect 12396 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12564 2752
rect 12244 2128 12564 2688
rect 13744 29408 14064 29424
rect 13744 29344 13752 29408
rect 13816 29344 13832 29408
rect 13896 29344 13912 29408
rect 13976 29344 13992 29408
rect 14056 29344 14064 29408
rect 13744 28320 14064 29344
rect 13744 28256 13752 28320
rect 13816 28256 13832 28320
rect 13896 28256 13912 28320
rect 13976 28256 13992 28320
rect 14056 28256 14064 28320
rect 13744 27232 14064 28256
rect 13744 27168 13752 27232
rect 13816 27168 13832 27232
rect 13896 27168 13912 27232
rect 13976 27168 13992 27232
rect 14056 27168 14064 27232
rect 13744 27046 14064 27168
rect 13744 26810 13786 27046
rect 14022 26810 14064 27046
rect 13744 26144 14064 26810
rect 13744 26080 13752 26144
rect 13816 26080 13832 26144
rect 13896 26080 13912 26144
rect 13976 26080 13992 26144
rect 14056 26080 14064 26144
rect 13744 25056 14064 26080
rect 13744 24992 13752 25056
rect 13816 24992 13832 25056
rect 13896 24992 13912 25056
rect 13976 24992 13992 25056
rect 14056 24992 14064 25056
rect 13744 24046 14064 24992
rect 13744 23968 13786 24046
rect 14022 23968 14064 24046
rect 13744 23904 13752 23968
rect 14056 23904 14064 23968
rect 13744 23810 13786 23904
rect 14022 23810 14064 23904
rect 13744 22880 14064 23810
rect 13744 22816 13752 22880
rect 13816 22816 13832 22880
rect 13896 22816 13912 22880
rect 13976 22816 13992 22880
rect 14056 22816 14064 22880
rect 13744 21792 14064 22816
rect 13744 21728 13752 21792
rect 13816 21728 13832 21792
rect 13896 21728 13912 21792
rect 13976 21728 13992 21792
rect 14056 21728 14064 21792
rect 13744 21046 14064 21728
rect 13744 20810 13786 21046
rect 14022 20810 14064 21046
rect 13744 20704 14064 20810
rect 13744 20640 13752 20704
rect 13816 20640 13832 20704
rect 13896 20640 13912 20704
rect 13976 20640 13992 20704
rect 14056 20640 14064 20704
rect 13744 19616 14064 20640
rect 13744 19552 13752 19616
rect 13816 19552 13832 19616
rect 13896 19552 13912 19616
rect 13976 19552 13992 19616
rect 14056 19552 14064 19616
rect 13744 18528 14064 19552
rect 13744 18464 13752 18528
rect 13816 18464 13832 18528
rect 13896 18464 13912 18528
rect 13976 18464 13992 18528
rect 14056 18464 14064 18528
rect 13744 18046 14064 18464
rect 13744 17810 13786 18046
rect 14022 17810 14064 18046
rect 13744 17440 14064 17810
rect 13744 17376 13752 17440
rect 13816 17376 13832 17440
rect 13896 17376 13912 17440
rect 13976 17376 13992 17440
rect 14056 17376 14064 17440
rect 13744 16352 14064 17376
rect 13744 16288 13752 16352
rect 13816 16288 13832 16352
rect 13896 16288 13912 16352
rect 13976 16288 13992 16352
rect 14056 16288 14064 16352
rect 13744 15264 14064 16288
rect 13744 15200 13752 15264
rect 13816 15200 13832 15264
rect 13896 15200 13912 15264
rect 13976 15200 13992 15264
rect 14056 15200 14064 15264
rect 13744 15046 14064 15200
rect 13744 14810 13786 15046
rect 14022 14810 14064 15046
rect 13744 14176 14064 14810
rect 13744 14112 13752 14176
rect 13816 14112 13832 14176
rect 13896 14112 13912 14176
rect 13976 14112 13992 14176
rect 14056 14112 14064 14176
rect 13744 13088 14064 14112
rect 13744 13024 13752 13088
rect 13816 13024 13832 13088
rect 13896 13024 13912 13088
rect 13976 13024 13992 13088
rect 14056 13024 14064 13088
rect 13744 12046 14064 13024
rect 13744 12000 13786 12046
rect 14022 12000 14064 12046
rect 13744 11936 13752 12000
rect 14056 11936 14064 12000
rect 13744 11810 13786 11936
rect 14022 11810 14064 11936
rect 13744 10912 14064 11810
rect 13744 10848 13752 10912
rect 13816 10848 13832 10912
rect 13896 10848 13912 10912
rect 13976 10848 13992 10912
rect 14056 10848 14064 10912
rect 13744 9824 14064 10848
rect 13744 9760 13752 9824
rect 13816 9760 13832 9824
rect 13896 9760 13912 9824
rect 13976 9760 13992 9824
rect 14056 9760 14064 9824
rect 13744 9046 14064 9760
rect 13744 8810 13786 9046
rect 14022 8810 14064 9046
rect 13744 8736 14064 8810
rect 13744 8672 13752 8736
rect 13816 8672 13832 8736
rect 13896 8672 13912 8736
rect 13976 8672 13992 8736
rect 14056 8672 14064 8736
rect 13744 7648 14064 8672
rect 13744 7584 13752 7648
rect 13816 7584 13832 7648
rect 13896 7584 13912 7648
rect 13976 7584 13992 7648
rect 14056 7584 14064 7648
rect 13744 6560 14064 7584
rect 13744 6496 13752 6560
rect 13816 6496 13832 6560
rect 13896 6496 13912 6560
rect 13976 6496 13992 6560
rect 14056 6496 14064 6560
rect 13744 6046 14064 6496
rect 13744 5810 13786 6046
rect 14022 5810 14064 6046
rect 13744 5472 14064 5810
rect 13744 5408 13752 5472
rect 13816 5408 13832 5472
rect 13896 5408 13912 5472
rect 13976 5408 13992 5472
rect 14056 5408 14064 5472
rect 13744 4384 14064 5408
rect 13744 4320 13752 4384
rect 13816 4320 13832 4384
rect 13896 4320 13912 4384
rect 13976 4320 13992 4384
rect 14056 4320 14064 4384
rect 13744 3296 14064 4320
rect 13744 3232 13752 3296
rect 13816 3232 13832 3296
rect 13896 3232 13912 3296
rect 13976 3232 13992 3296
rect 14056 3232 14064 3296
rect 13744 3046 14064 3232
rect 13744 2810 13786 3046
rect 14022 2810 14064 3046
rect 13744 2208 14064 2810
rect 13744 2144 13752 2208
rect 13816 2144 13832 2208
rect 13896 2144 13912 2208
rect 13976 2144 13992 2208
rect 14056 2144 14064 2208
rect 13744 2128 14064 2144
rect 15244 28864 15564 29424
rect 15244 28800 15252 28864
rect 15316 28800 15332 28864
rect 15396 28800 15412 28864
rect 15476 28800 15492 28864
rect 15556 28800 15564 28864
rect 15244 28546 15564 28800
rect 15244 28310 15286 28546
rect 15522 28310 15564 28546
rect 15244 27776 15564 28310
rect 15244 27712 15252 27776
rect 15316 27712 15332 27776
rect 15396 27712 15412 27776
rect 15476 27712 15492 27776
rect 15556 27712 15564 27776
rect 15244 26688 15564 27712
rect 15244 26624 15252 26688
rect 15316 26624 15332 26688
rect 15396 26624 15412 26688
rect 15476 26624 15492 26688
rect 15556 26624 15564 26688
rect 15244 25600 15564 26624
rect 15244 25536 15252 25600
rect 15316 25546 15332 25600
rect 15396 25546 15412 25600
rect 15476 25546 15492 25600
rect 15556 25536 15564 25600
rect 15244 25310 15286 25536
rect 15522 25310 15564 25536
rect 15244 24512 15564 25310
rect 15244 24448 15252 24512
rect 15316 24448 15332 24512
rect 15396 24448 15412 24512
rect 15476 24448 15492 24512
rect 15556 24448 15564 24512
rect 15244 23424 15564 24448
rect 15244 23360 15252 23424
rect 15316 23360 15332 23424
rect 15396 23360 15412 23424
rect 15476 23360 15492 23424
rect 15556 23360 15564 23424
rect 15244 22546 15564 23360
rect 15244 22336 15286 22546
rect 15522 22336 15564 22546
rect 15244 22272 15252 22336
rect 15316 22272 15332 22310
rect 15396 22272 15412 22310
rect 15476 22272 15492 22310
rect 15556 22272 15564 22336
rect 15244 21248 15564 22272
rect 15244 21184 15252 21248
rect 15316 21184 15332 21248
rect 15396 21184 15412 21248
rect 15476 21184 15492 21248
rect 15556 21184 15564 21248
rect 15244 20160 15564 21184
rect 15244 20096 15252 20160
rect 15316 20096 15332 20160
rect 15396 20096 15412 20160
rect 15476 20096 15492 20160
rect 15556 20096 15564 20160
rect 15244 19546 15564 20096
rect 15244 19310 15286 19546
rect 15522 19310 15564 19546
rect 15244 19072 15564 19310
rect 15244 19008 15252 19072
rect 15316 19008 15332 19072
rect 15396 19008 15412 19072
rect 15476 19008 15492 19072
rect 15556 19008 15564 19072
rect 15244 17984 15564 19008
rect 15244 17920 15252 17984
rect 15316 17920 15332 17984
rect 15396 17920 15412 17984
rect 15476 17920 15492 17984
rect 15556 17920 15564 17984
rect 15244 16896 15564 17920
rect 15244 16832 15252 16896
rect 15316 16832 15332 16896
rect 15396 16832 15412 16896
rect 15476 16832 15492 16896
rect 15556 16832 15564 16896
rect 15244 16546 15564 16832
rect 15244 16310 15286 16546
rect 15522 16310 15564 16546
rect 15244 15808 15564 16310
rect 15244 15744 15252 15808
rect 15316 15744 15332 15808
rect 15396 15744 15412 15808
rect 15476 15744 15492 15808
rect 15556 15744 15564 15808
rect 15244 14720 15564 15744
rect 15244 14656 15252 14720
rect 15316 14656 15332 14720
rect 15396 14656 15412 14720
rect 15476 14656 15492 14720
rect 15556 14656 15564 14720
rect 15244 13632 15564 14656
rect 15244 13568 15252 13632
rect 15316 13568 15332 13632
rect 15396 13568 15412 13632
rect 15476 13568 15492 13632
rect 15556 13568 15564 13632
rect 15244 13546 15564 13568
rect 15244 13310 15286 13546
rect 15522 13310 15564 13546
rect 15244 12544 15564 13310
rect 15244 12480 15252 12544
rect 15316 12480 15332 12544
rect 15396 12480 15412 12544
rect 15476 12480 15492 12544
rect 15556 12480 15564 12544
rect 15244 11456 15564 12480
rect 15244 11392 15252 11456
rect 15316 11392 15332 11456
rect 15396 11392 15412 11456
rect 15476 11392 15492 11456
rect 15556 11392 15564 11456
rect 15244 10546 15564 11392
rect 15244 10368 15286 10546
rect 15522 10368 15564 10546
rect 15244 10304 15252 10368
rect 15316 10304 15332 10310
rect 15396 10304 15412 10310
rect 15476 10304 15492 10310
rect 15556 10304 15564 10368
rect 15244 9280 15564 10304
rect 15244 9216 15252 9280
rect 15316 9216 15332 9280
rect 15396 9216 15412 9280
rect 15476 9216 15492 9280
rect 15556 9216 15564 9280
rect 15244 8192 15564 9216
rect 15244 8128 15252 8192
rect 15316 8128 15332 8192
rect 15396 8128 15412 8192
rect 15476 8128 15492 8192
rect 15556 8128 15564 8192
rect 15244 7546 15564 8128
rect 15244 7310 15286 7546
rect 15522 7310 15564 7546
rect 15244 7104 15564 7310
rect 15244 7040 15252 7104
rect 15316 7040 15332 7104
rect 15396 7040 15412 7104
rect 15476 7040 15492 7104
rect 15556 7040 15564 7104
rect 15244 6016 15564 7040
rect 15244 5952 15252 6016
rect 15316 5952 15332 6016
rect 15396 5952 15412 6016
rect 15476 5952 15492 6016
rect 15556 5952 15564 6016
rect 15244 4928 15564 5952
rect 15244 4864 15252 4928
rect 15316 4864 15332 4928
rect 15396 4864 15412 4928
rect 15476 4864 15492 4928
rect 15556 4864 15564 4928
rect 15244 4546 15564 4864
rect 15244 4310 15286 4546
rect 15522 4310 15564 4546
rect 15244 3840 15564 4310
rect 15244 3776 15252 3840
rect 15316 3776 15332 3840
rect 15396 3776 15412 3840
rect 15476 3776 15492 3840
rect 15556 3776 15564 3840
rect 15244 2752 15564 3776
rect 15244 2688 15252 2752
rect 15316 2688 15332 2752
rect 15396 2688 15412 2752
rect 15476 2688 15492 2752
rect 15556 2688 15564 2752
rect 15244 2128 15564 2688
rect 16744 29408 17064 29424
rect 16744 29344 16752 29408
rect 16816 29344 16832 29408
rect 16896 29344 16912 29408
rect 16976 29344 16992 29408
rect 17056 29344 17064 29408
rect 16744 28320 17064 29344
rect 16744 28256 16752 28320
rect 16816 28256 16832 28320
rect 16896 28256 16912 28320
rect 16976 28256 16992 28320
rect 17056 28256 17064 28320
rect 16744 27232 17064 28256
rect 16744 27168 16752 27232
rect 16816 27168 16832 27232
rect 16896 27168 16912 27232
rect 16976 27168 16992 27232
rect 17056 27168 17064 27232
rect 16744 27046 17064 27168
rect 16744 26810 16786 27046
rect 17022 26810 17064 27046
rect 16744 26144 17064 26810
rect 16744 26080 16752 26144
rect 16816 26080 16832 26144
rect 16896 26080 16912 26144
rect 16976 26080 16992 26144
rect 17056 26080 17064 26144
rect 16744 25056 17064 26080
rect 16744 24992 16752 25056
rect 16816 24992 16832 25056
rect 16896 24992 16912 25056
rect 16976 24992 16992 25056
rect 17056 24992 17064 25056
rect 16744 24046 17064 24992
rect 16744 23968 16786 24046
rect 17022 23968 17064 24046
rect 16744 23904 16752 23968
rect 17056 23904 17064 23968
rect 16744 23810 16786 23904
rect 17022 23810 17064 23904
rect 16744 22880 17064 23810
rect 16744 22816 16752 22880
rect 16816 22816 16832 22880
rect 16896 22816 16912 22880
rect 16976 22816 16992 22880
rect 17056 22816 17064 22880
rect 16744 21792 17064 22816
rect 16744 21728 16752 21792
rect 16816 21728 16832 21792
rect 16896 21728 16912 21792
rect 16976 21728 16992 21792
rect 17056 21728 17064 21792
rect 16744 21046 17064 21728
rect 16744 20810 16786 21046
rect 17022 20810 17064 21046
rect 16744 20704 17064 20810
rect 16744 20640 16752 20704
rect 16816 20640 16832 20704
rect 16896 20640 16912 20704
rect 16976 20640 16992 20704
rect 17056 20640 17064 20704
rect 16744 19616 17064 20640
rect 16744 19552 16752 19616
rect 16816 19552 16832 19616
rect 16896 19552 16912 19616
rect 16976 19552 16992 19616
rect 17056 19552 17064 19616
rect 16744 18528 17064 19552
rect 16744 18464 16752 18528
rect 16816 18464 16832 18528
rect 16896 18464 16912 18528
rect 16976 18464 16992 18528
rect 17056 18464 17064 18528
rect 16744 18046 17064 18464
rect 16744 17810 16786 18046
rect 17022 17810 17064 18046
rect 16744 17440 17064 17810
rect 16744 17376 16752 17440
rect 16816 17376 16832 17440
rect 16896 17376 16912 17440
rect 16976 17376 16992 17440
rect 17056 17376 17064 17440
rect 16744 16352 17064 17376
rect 16744 16288 16752 16352
rect 16816 16288 16832 16352
rect 16896 16288 16912 16352
rect 16976 16288 16992 16352
rect 17056 16288 17064 16352
rect 16744 15264 17064 16288
rect 16744 15200 16752 15264
rect 16816 15200 16832 15264
rect 16896 15200 16912 15264
rect 16976 15200 16992 15264
rect 17056 15200 17064 15264
rect 16744 15046 17064 15200
rect 16744 14810 16786 15046
rect 17022 14810 17064 15046
rect 16744 14176 17064 14810
rect 16744 14112 16752 14176
rect 16816 14112 16832 14176
rect 16896 14112 16912 14176
rect 16976 14112 16992 14176
rect 17056 14112 17064 14176
rect 16744 13088 17064 14112
rect 16744 13024 16752 13088
rect 16816 13024 16832 13088
rect 16896 13024 16912 13088
rect 16976 13024 16992 13088
rect 17056 13024 17064 13088
rect 16744 12046 17064 13024
rect 16744 12000 16786 12046
rect 17022 12000 17064 12046
rect 16744 11936 16752 12000
rect 17056 11936 17064 12000
rect 16744 11810 16786 11936
rect 17022 11810 17064 11936
rect 16744 10912 17064 11810
rect 16744 10848 16752 10912
rect 16816 10848 16832 10912
rect 16896 10848 16912 10912
rect 16976 10848 16992 10912
rect 17056 10848 17064 10912
rect 16744 9824 17064 10848
rect 16744 9760 16752 9824
rect 16816 9760 16832 9824
rect 16896 9760 16912 9824
rect 16976 9760 16992 9824
rect 17056 9760 17064 9824
rect 16744 9046 17064 9760
rect 16744 8810 16786 9046
rect 17022 8810 17064 9046
rect 16744 8736 17064 8810
rect 16744 8672 16752 8736
rect 16816 8672 16832 8736
rect 16896 8672 16912 8736
rect 16976 8672 16992 8736
rect 17056 8672 17064 8736
rect 16744 7648 17064 8672
rect 16744 7584 16752 7648
rect 16816 7584 16832 7648
rect 16896 7584 16912 7648
rect 16976 7584 16992 7648
rect 17056 7584 17064 7648
rect 16744 6560 17064 7584
rect 16744 6496 16752 6560
rect 16816 6496 16832 6560
rect 16896 6496 16912 6560
rect 16976 6496 16992 6560
rect 17056 6496 17064 6560
rect 16744 6046 17064 6496
rect 16744 5810 16786 6046
rect 17022 5810 17064 6046
rect 16744 5472 17064 5810
rect 16744 5408 16752 5472
rect 16816 5408 16832 5472
rect 16896 5408 16912 5472
rect 16976 5408 16992 5472
rect 17056 5408 17064 5472
rect 16744 4384 17064 5408
rect 16744 4320 16752 4384
rect 16816 4320 16832 4384
rect 16896 4320 16912 4384
rect 16976 4320 16992 4384
rect 17056 4320 17064 4384
rect 16744 3296 17064 4320
rect 16744 3232 16752 3296
rect 16816 3232 16832 3296
rect 16896 3232 16912 3296
rect 16976 3232 16992 3296
rect 17056 3232 17064 3296
rect 16744 3046 17064 3232
rect 16744 2810 16786 3046
rect 17022 2810 17064 3046
rect 16744 2208 17064 2810
rect 16744 2144 16752 2208
rect 16816 2144 16832 2208
rect 16896 2144 16912 2208
rect 16976 2144 16992 2208
rect 17056 2144 17064 2208
rect 16744 2128 17064 2144
rect 18244 28864 18564 29424
rect 18244 28800 18252 28864
rect 18316 28800 18332 28864
rect 18396 28800 18412 28864
rect 18476 28800 18492 28864
rect 18556 28800 18564 28864
rect 18244 28546 18564 28800
rect 18244 28310 18286 28546
rect 18522 28310 18564 28546
rect 18244 27776 18564 28310
rect 18244 27712 18252 27776
rect 18316 27712 18332 27776
rect 18396 27712 18412 27776
rect 18476 27712 18492 27776
rect 18556 27712 18564 27776
rect 18244 26688 18564 27712
rect 18244 26624 18252 26688
rect 18316 26624 18332 26688
rect 18396 26624 18412 26688
rect 18476 26624 18492 26688
rect 18556 26624 18564 26688
rect 18244 25600 18564 26624
rect 18244 25536 18252 25600
rect 18316 25546 18332 25600
rect 18396 25546 18412 25600
rect 18476 25546 18492 25600
rect 18556 25536 18564 25600
rect 18244 25310 18286 25536
rect 18522 25310 18564 25536
rect 18244 24512 18564 25310
rect 18244 24448 18252 24512
rect 18316 24448 18332 24512
rect 18396 24448 18412 24512
rect 18476 24448 18492 24512
rect 18556 24448 18564 24512
rect 18244 23424 18564 24448
rect 18244 23360 18252 23424
rect 18316 23360 18332 23424
rect 18396 23360 18412 23424
rect 18476 23360 18492 23424
rect 18556 23360 18564 23424
rect 18244 22546 18564 23360
rect 18244 22336 18286 22546
rect 18522 22336 18564 22546
rect 18244 22272 18252 22336
rect 18316 22272 18332 22310
rect 18396 22272 18412 22310
rect 18476 22272 18492 22310
rect 18556 22272 18564 22336
rect 18244 21248 18564 22272
rect 18244 21184 18252 21248
rect 18316 21184 18332 21248
rect 18396 21184 18412 21248
rect 18476 21184 18492 21248
rect 18556 21184 18564 21248
rect 18244 20160 18564 21184
rect 18244 20096 18252 20160
rect 18316 20096 18332 20160
rect 18396 20096 18412 20160
rect 18476 20096 18492 20160
rect 18556 20096 18564 20160
rect 18244 19546 18564 20096
rect 18244 19310 18286 19546
rect 18522 19310 18564 19546
rect 18244 19072 18564 19310
rect 18244 19008 18252 19072
rect 18316 19008 18332 19072
rect 18396 19008 18412 19072
rect 18476 19008 18492 19072
rect 18556 19008 18564 19072
rect 18244 17984 18564 19008
rect 18244 17920 18252 17984
rect 18316 17920 18332 17984
rect 18396 17920 18412 17984
rect 18476 17920 18492 17984
rect 18556 17920 18564 17984
rect 18244 16896 18564 17920
rect 18244 16832 18252 16896
rect 18316 16832 18332 16896
rect 18396 16832 18412 16896
rect 18476 16832 18492 16896
rect 18556 16832 18564 16896
rect 18244 16546 18564 16832
rect 18244 16310 18286 16546
rect 18522 16310 18564 16546
rect 18244 15808 18564 16310
rect 18244 15744 18252 15808
rect 18316 15744 18332 15808
rect 18396 15744 18412 15808
rect 18476 15744 18492 15808
rect 18556 15744 18564 15808
rect 18244 14720 18564 15744
rect 18244 14656 18252 14720
rect 18316 14656 18332 14720
rect 18396 14656 18412 14720
rect 18476 14656 18492 14720
rect 18556 14656 18564 14720
rect 18244 13632 18564 14656
rect 19744 29408 20064 29424
rect 19744 29344 19752 29408
rect 19816 29344 19832 29408
rect 19896 29344 19912 29408
rect 19976 29344 19992 29408
rect 20056 29344 20064 29408
rect 19744 28320 20064 29344
rect 19744 28256 19752 28320
rect 19816 28256 19832 28320
rect 19896 28256 19912 28320
rect 19976 28256 19992 28320
rect 20056 28256 20064 28320
rect 19744 27232 20064 28256
rect 19744 27168 19752 27232
rect 19816 27168 19832 27232
rect 19896 27168 19912 27232
rect 19976 27168 19992 27232
rect 20056 27168 20064 27232
rect 19744 27046 20064 27168
rect 19744 26810 19786 27046
rect 20022 26810 20064 27046
rect 19744 26144 20064 26810
rect 19744 26080 19752 26144
rect 19816 26080 19832 26144
rect 19896 26080 19912 26144
rect 19976 26080 19992 26144
rect 20056 26080 20064 26144
rect 19744 25056 20064 26080
rect 19744 24992 19752 25056
rect 19816 24992 19832 25056
rect 19896 24992 19912 25056
rect 19976 24992 19992 25056
rect 20056 24992 20064 25056
rect 19744 24046 20064 24992
rect 19744 23968 19786 24046
rect 20022 23968 20064 24046
rect 19744 23904 19752 23968
rect 20056 23904 20064 23968
rect 19744 23810 19786 23904
rect 20022 23810 20064 23904
rect 19744 22880 20064 23810
rect 19744 22816 19752 22880
rect 19816 22816 19832 22880
rect 19896 22816 19912 22880
rect 19976 22816 19992 22880
rect 20056 22816 20064 22880
rect 19744 21792 20064 22816
rect 19744 21728 19752 21792
rect 19816 21728 19832 21792
rect 19896 21728 19912 21792
rect 19976 21728 19992 21792
rect 20056 21728 20064 21792
rect 19744 21046 20064 21728
rect 19744 20810 19786 21046
rect 20022 20810 20064 21046
rect 19744 20704 20064 20810
rect 19744 20640 19752 20704
rect 19816 20640 19832 20704
rect 19896 20640 19912 20704
rect 19976 20640 19992 20704
rect 20056 20640 20064 20704
rect 19744 19616 20064 20640
rect 19744 19552 19752 19616
rect 19816 19552 19832 19616
rect 19896 19552 19912 19616
rect 19976 19552 19992 19616
rect 20056 19552 20064 19616
rect 19744 18528 20064 19552
rect 19744 18464 19752 18528
rect 19816 18464 19832 18528
rect 19896 18464 19912 18528
rect 19976 18464 19992 18528
rect 20056 18464 20064 18528
rect 19744 18046 20064 18464
rect 19744 17810 19786 18046
rect 20022 17810 20064 18046
rect 19744 17440 20064 17810
rect 19744 17376 19752 17440
rect 19816 17376 19832 17440
rect 19896 17376 19912 17440
rect 19976 17376 19992 17440
rect 20056 17376 20064 17440
rect 19744 16352 20064 17376
rect 19744 16288 19752 16352
rect 19816 16288 19832 16352
rect 19896 16288 19912 16352
rect 19976 16288 19992 16352
rect 20056 16288 20064 16352
rect 19744 15264 20064 16288
rect 19744 15200 19752 15264
rect 19816 15200 19832 15264
rect 19896 15200 19912 15264
rect 19976 15200 19992 15264
rect 20056 15200 20064 15264
rect 19744 15046 20064 15200
rect 19744 14810 19786 15046
rect 20022 14810 20064 15046
rect 19379 14516 19445 14517
rect 19379 14452 19380 14516
rect 19444 14452 19445 14516
rect 19379 14451 19445 14452
rect 18244 13568 18252 13632
rect 18316 13568 18332 13632
rect 18396 13568 18412 13632
rect 18476 13568 18492 13632
rect 18556 13568 18564 13632
rect 18244 13546 18564 13568
rect 18244 13310 18286 13546
rect 18522 13310 18564 13546
rect 18244 12544 18564 13310
rect 18244 12480 18252 12544
rect 18316 12480 18332 12544
rect 18396 12480 18412 12544
rect 18476 12480 18492 12544
rect 18556 12480 18564 12544
rect 18244 11456 18564 12480
rect 18244 11392 18252 11456
rect 18316 11392 18332 11456
rect 18396 11392 18412 11456
rect 18476 11392 18492 11456
rect 18556 11392 18564 11456
rect 18244 10546 18564 11392
rect 18244 10368 18286 10546
rect 18522 10368 18564 10546
rect 18244 10304 18252 10368
rect 18316 10304 18332 10310
rect 18396 10304 18412 10310
rect 18476 10304 18492 10310
rect 18556 10304 18564 10368
rect 18244 9280 18564 10304
rect 19382 10029 19442 14451
rect 19744 14176 20064 14810
rect 19744 14112 19752 14176
rect 19816 14112 19832 14176
rect 19896 14112 19912 14176
rect 19976 14112 19992 14176
rect 20056 14112 20064 14176
rect 19744 13088 20064 14112
rect 19744 13024 19752 13088
rect 19816 13024 19832 13088
rect 19896 13024 19912 13088
rect 19976 13024 19992 13088
rect 20056 13024 20064 13088
rect 19744 12046 20064 13024
rect 19744 12000 19786 12046
rect 20022 12000 20064 12046
rect 19744 11936 19752 12000
rect 20056 11936 20064 12000
rect 19744 11810 19786 11936
rect 20022 11810 20064 11936
rect 19744 10912 20064 11810
rect 19744 10848 19752 10912
rect 19816 10848 19832 10912
rect 19896 10848 19912 10912
rect 19976 10848 19992 10912
rect 20056 10848 20064 10912
rect 19379 10028 19445 10029
rect 19379 9964 19380 10028
rect 19444 9964 19445 10028
rect 19379 9963 19445 9964
rect 18244 9216 18252 9280
rect 18316 9216 18332 9280
rect 18396 9216 18412 9280
rect 18476 9216 18492 9280
rect 18556 9216 18564 9280
rect 18244 8192 18564 9216
rect 18244 8128 18252 8192
rect 18316 8128 18332 8192
rect 18396 8128 18412 8192
rect 18476 8128 18492 8192
rect 18556 8128 18564 8192
rect 18244 7546 18564 8128
rect 18244 7310 18286 7546
rect 18522 7310 18564 7546
rect 18244 7104 18564 7310
rect 18244 7040 18252 7104
rect 18316 7040 18332 7104
rect 18396 7040 18412 7104
rect 18476 7040 18492 7104
rect 18556 7040 18564 7104
rect 18244 6016 18564 7040
rect 18244 5952 18252 6016
rect 18316 5952 18332 6016
rect 18396 5952 18412 6016
rect 18476 5952 18492 6016
rect 18556 5952 18564 6016
rect 18244 4928 18564 5952
rect 18244 4864 18252 4928
rect 18316 4864 18332 4928
rect 18396 4864 18412 4928
rect 18476 4864 18492 4928
rect 18556 4864 18564 4928
rect 18244 4546 18564 4864
rect 18244 4310 18286 4546
rect 18522 4310 18564 4546
rect 18244 3840 18564 4310
rect 18244 3776 18252 3840
rect 18316 3776 18332 3840
rect 18396 3776 18412 3840
rect 18476 3776 18492 3840
rect 18556 3776 18564 3840
rect 18244 2752 18564 3776
rect 18244 2688 18252 2752
rect 18316 2688 18332 2752
rect 18396 2688 18412 2752
rect 18476 2688 18492 2752
rect 18556 2688 18564 2752
rect 18244 2128 18564 2688
rect 19744 9824 20064 10848
rect 19744 9760 19752 9824
rect 19816 9760 19832 9824
rect 19896 9760 19912 9824
rect 19976 9760 19992 9824
rect 20056 9760 20064 9824
rect 19744 9046 20064 9760
rect 19744 8810 19786 9046
rect 20022 8810 20064 9046
rect 19744 8736 20064 8810
rect 19744 8672 19752 8736
rect 19816 8672 19832 8736
rect 19896 8672 19912 8736
rect 19976 8672 19992 8736
rect 20056 8672 20064 8736
rect 19744 7648 20064 8672
rect 19744 7584 19752 7648
rect 19816 7584 19832 7648
rect 19896 7584 19912 7648
rect 19976 7584 19992 7648
rect 20056 7584 20064 7648
rect 19744 6560 20064 7584
rect 19744 6496 19752 6560
rect 19816 6496 19832 6560
rect 19896 6496 19912 6560
rect 19976 6496 19992 6560
rect 20056 6496 20064 6560
rect 19744 6046 20064 6496
rect 19744 5810 19786 6046
rect 20022 5810 20064 6046
rect 19744 5472 20064 5810
rect 19744 5408 19752 5472
rect 19816 5408 19832 5472
rect 19896 5408 19912 5472
rect 19976 5408 19992 5472
rect 20056 5408 20064 5472
rect 19744 4384 20064 5408
rect 19744 4320 19752 4384
rect 19816 4320 19832 4384
rect 19896 4320 19912 4384
rect 19976 4320 19992 4384
rect 20056 4320 20064 4384
rect 19744 3296 20064 4320
rect 19744 3232 19752 3296
rect 19816 3232 19832 3296
rect 19896 3232 19912 3296
rect 19976 3232 19992 3296
rect 20056 3232 20064 3296
rect 19744 3046 20064 3232
rect 19744 2810 19786 3046
rect 20022 2810 20064 3046
rect 19744 2208 20064 2810
rect 19744 2144 19752 2208
rect 19816 2144 19832 2208
rect 19896 2144 19912 2208
rect 19976 2144 19992 2208
rect 20056 2144 20064 2208
rect 19744 2128 20064 2144
rect 21244 28864 21564 29424
rect 21244 28800 21252 28864
rect 21316 28800 21332 28864
rect 21396 28800 21412 28864
rect 21476 28800 21492 28864
rect 21556 28800 21564 28864
rect 21244 28546 21564 28800
rect 21244 28310 21286 28546
rect 21522 28310 21564 28546
rect 21244 27776 21564 28310
rect 21244 27712 21252 27776
rect 21316 27712 21332 27776
rect 21396 27712 21412 27776
rect 21476 27712 21492 27776
rect 21556 27712 21564 27776
rect 21244 26688 21564 27712
rect 21244 26624 21252 26688
rect 21316 26624 21332 26688
rect 21396 26624 21412 26688
rect 21476 26624 21492 26688
rect 21556 26624 21564 26688
rect 21244 25600 21564 26624
rect 21244 25536 21252 25600
rect 21316 25546 21332 25600
rect 21396 25546 21412 25600
rect 21476 25546 21492 25600
rect 21556 25536 21564 25600
rect 21244 25310 21286 25536
rect 21522 25310 21564 25536
rect 21244 24512 21564 25310
rect 21244 24448 21252 24512
rect 21316 24448 21332 24512
rect 21396 24448 21412 24512
rect 21476 24448 21492 24512
rect 21556 24448 21564 24512
rect 21244 23424 21564 24448
rect 21244 23360 21252 23424
rect 21316 23360 21332 23424
rect 21396 23360 21412 23424
rect 21476 23360 21492 23424
rect 21556 23360 21564 23424
rect 21244 22546 21564 23360
rect 21244 22336 21286 22546
rect 21522 22336 21564 22546
rect 21244 22272 21252 22336
rect 21316 22272 21332 22310
rect 21396 22272 21412 22310
rect 21476 22272 21492 22310
rect 21556 22272 21564 22336
rect 21244 21248 21564 22272
rect 21244 21184 21252 21248
rect 21316 21184 21332 21248
rect 21396 21184 21412 21248
rect 21476 21184 21492 21248
rect 21556 21184 21564 21248
rect 21244 20160 21564 21184
rect 21244 20096 21252 20160
rect 21316 20096 21332 20160
rect 21396 20096 21412 20160
rect 21476 20096 21492 20160
rect 21556 20096 21564 20160
rect 21244 19546 21564 20096
rect 21244 19310 21286 19546
rect 21522 19310 21564 19546
rect 21244 19072 21564 19310
rect 21244 19008 21252 19072
rect 21316 19008 21332 19072
rect 21396 19008 21412 19072
rect 21476 19008 21492 19072
rect 21556 19008 21564 19072
rect 21244 17984 21564 19008
rect 21244 17920 21252 17984
rect 21316 17920 21332 17984
rect 21396 17920 21412 17984
rect 21476 17920 21492 17984
rect 21556 17920 21564 17984
rect 21244 16896 21564 17920
rect 21244 16832 21252 16896
rect 21316 16832 21332 16896
rect 21396 16832 21412 16896
rect 21476 16832 21492 16896
rect 21556 16832 21564 16896
rect 21244 16546 21564 16832
rect 21244 16310 21286 16546
rect 21522 16310 21564 16546
rect 21244 15808 21564 16310
rect 21244 15744 21252 15808
rect 21316 15744 21332 15808
rect 21396 15744 21412 15808
rect 21476 15744 21492 15808
rect 21556 15744 21564 15808
rect 21244 14720 21564 15744
rect 21244 14656 21252 14720
rect 21316 14656 21332 14720
rect 21396 14656 21412 14720
rect 21476 14656 21492 14720
rect 21556 14656 21564 14720
rect 21244 13632 21564 14656
rect 21244 13568 21252 13632
rect 21316 13568 21332 13632
rect 21396 13568 21412 13632
rect 21476 13568 21492 13632
rect 21556 13568 21564 13632
rect 21244 13546 21564 13568
rect 21244 13310 21286 13546
rect 21522 13310 21564 13546
rect 21244 12544 21564 13310
rect 21244 12480 21252 12544
rect 21316 12480 21332 12544
rect 21396 12480 21412 12544
rect 21476 12480 21492 12544
rect 21556 12480 21564 12544
rect 21244 11456 21564 12480
rect 21244 11392 21252 11456
rect 21316 11392 21332 11456
rect 21396 11392 21412 11456
rect 21476 11392 21492 11456
rect 21556 11392 21564 11456
rect 21244 10546 21564 11392
rect 21244 10368 21286 10546
rect 21522 10368 21564 10546
rect 21244 10304 21252 10368
rect 21316 10304 21332 10310
rect 21396 10304 21412 10310
rect 21476 10304 21492 10310
rect 21556 10304 21564 10368
rect 21244 9280 21564 10304
rect 21244 9216 21252 9280
rect 21316 9216 21332 9280
rect 21396 9216 21412 9280
rect 21476 9216 21492 9280
rect 21556 9216 21564 9280
rect 21244 8192 21564 9216
rect 21244 8128 21252 8192
rect 21316 8128 21332 8192
rect 21396 8128 21412 8192
rect 21476 8128 21492 8192
rect 21556 8128 21564 8192
rect 21244 7546 21564 8128
rect 21244 7310 21286 7546
rect 21522 7310 21564 7546
rect 21244 7104 21564 7310
rect 21244 7040 21252 7104
rect 21316 7040 21332 7104
rect 21396 7040 21412 7104
rect 21476 7040 21492 7104
rect 21556 7040 21564 7104
rect 21244 6016 21564 7040
rect 21244 5952 21252 6016
rect 21316 5952 21332 6016
rect 21396 5952 21412 6016
rect 21476 5952 21492 6016
rect 21556 5952 21564 6016
rect 21244 4928 21564 5952
rect 21244 4864 21252 4928
rect 21316 4864 21332 4928
rect 21396 4864 21412 4928
rect 21476 4864 21492 4928
rect 21556 4864 21564 4928
rect 21244 4546 21564 4864
rect 21244 4310 21286 4546
rect 21522 4310 21564 4546
rect 21244 3840 21564 4310
rect 21244 3776 21252 3840
rect 21316 3776 21332 3840
rect 21396 3776 21412 3840
rect 21476 3776 21492 3840
rect 21556 3776 21564 3840
rect 21244 2752 21564 3776
rect 21244 2688 21252 2752
rect 21316 2688 21332 2752
rect 21396 2688 21412 2752
rect 21476 2688 21492 2752
rect 21556 2688 21564 2752
rect 21244 2128 21564 2688
rect 22744 29408 23064 29424
rect 22744 29344 22752 29408
rect 22816 29344 22832 29408
rect 22896 29344 22912 29408
rect 22976 29344 22992 29408
rect 23056 29344 23064 29408
rect 22744 28320 23064 29344
rect 22744 28256 22752 28320
rect 22816 28256 22832 28320
rect 22896 28256 22912 28320
rect 22976 28256 22992 28320
rect 23056 28256 23064 28320
rect 22744 27232 23064 28256
rect 22744 27168 22752 27232
rect 22816 27168 22832 27232
rect 22896 27168 22912 27232
rect 22976 27168 22992 27232
rect 23056 27168 23064 27232
rect 22744 27046 23064 27168
rect 22744 26810 22786 27046
rect 23022 26810 23064 27046
rect 22744 26144 23064 26810
rect 22744 26080 22752 26144
rect 22816 26080 22832 26144
rect 22896 26080 22912 26144
rect 22976 26080 22992 26144
rect 23056 26080 23064 26144
rect 22744 25056 23064 26080
rect 22744 24992 22752 25056
rect 22816 24992 22832 25056
rect 22896 24992 22912 25056
rect 22976 24992 22992 25056
rect 23056 24992 23064 25056
rect 22744 24046 23064 24992
rect 22744 23968 22786 24046
rect 23022 23968 23064 24046
rect 22744 23904 22752 23968
rect 23056 23904 23064 23968
rect 22744 23810 22786 23904
rect 23022 23810 23064 23904
rect 22744 22880 23064 23810
rect 22744 22816 22752 22880
rect 22816 22816 22832 22880
rect 22896 22816 22912 22880
rect 22976 22816 22992 22880
rect 23056 22816 23064 22880
rect 22744 21792 23064 22816
rect 22744 21728 22752 21792
rect 22816 21728 22832 21792
rect 22896 21728 22912 21792
rect 22976 21728 22992 21792
rect 23056 21728 23064 21792
rect 22744 21046 23064 21728
rect 22744 20810 22786 21046
rect 23022 20810 23064 21046
rect 22744 20704 23064 20810
rect 22744 20640 22752 20704
rect 22816 20640 22832 20704
rect 22896 20640 22912 20704
rect 22976 20640 22992 20704
rect 23056 20640 23064 20704
rect 22744 19616 23064 20640
rect 22744 19552 22752 19616
rect 22816 19552 22832 19616
rect 22896 19552 22912 19616
rect 22976 19552 22992 19616
rect 23056 19552 23064 19616
rect 22744 18528 23064 19552
rect 22744 18464 22752 18528
rect 22816 18464 22832 18528
rect 22896 18464 22912 18528
rect 22976 18464 22992 18528
rect 23056 18464 23064 18528
rect 22744 18046 23064 18464
rect 22744 17810 22786 18046
rect 23022 17810 23064 18046
rect 22744 17440 23064 17810
rect 22744 17376 22752 17440
rect 22816 17376 22832 17440
rect 22896 17376 22912 17440
rect 22976 17376 22992 17440
rect 23056 17376 23064 17440
rect 22744 16352 23064 17376
rect 22744 16288 22752 16352
rect 22816 16288 22832 16352
rect 22896 16288 22912 16352
rect 22976 16288 22992 16352
rect 23056 16288 23064 16352
rect 22744 15264 23064 16288
rect 22744 15200 22752 15264
rect 22816 15200 22832 15264
rect 22896 15200 22912 15264
rect 22976 15200 22992 15264
rect 23056 15200 23064 15264
rect 22744 15046 23064 15200
rect 22744 14810 22786 15046
rect 23022 14810 23064 15046
rect 22744 14176 23064 14810
rect 22744 14112 22752 14176
rect 22816 14112 22832 14176
rect 22896 14112 22912 14176
rect 22976 14112 22992 14176
rect 23056 14112 23064 14176
rect 22744 13088 23064 14112
rect 22744 13024 22752 13088
rect 22816 13024 22832 13088
rect 22896 13024 22912 13088
rect 22976 13024 22992 13088
rect 23056 13024 23064 13088
rect 22744 12046 23064 13024
rect 22744 12000 22786 12046
rect 23022 12000 23064 12046
rect 22744 11936 22752 12000
rect 23056 11936 23064 12000
rect 22744 11810 22786 11936
rect 23022 11810 23064 11936
rect 22744 10912 23064 11810
rect 22744 10848 22752 10912
rect 22816 10848 22832 10912
rect 22896 10848 22912 10912
rect 22976 10848 22992 10912
rect 23056 10848 23064 10912
rect 22744 9824 23064 10848
rect 22744 9760 22752 9824
rect 22816 9760 22832 9824
rect 22896 9760 22912 9824
rect 22976 9760 22992 9824
rect 23056 9760 23064 9824
rect 22744 9046 23064 9760
rect 22744 8810 22786 9046
rect 23022 8810 23064 9046
rect 22744 8736 23064 8810
rect 22744 8672 22752 8736
rect 22816 8672 22832 8736
rect 22896 8672 22912 8736
rect 22976 8672 22992 8736
rect 23056 8672 23064 8736
rect 22744 7648 23064 8672
rect 22744 7584 22752 7648
rect 22816 7584 22832 7648
rect 22896 7584 22912 7648
rect 22976 7584 22992 7648
rect 23056 7584 23064 7648
rect 22744 6560 23064 7584
rect 22744 6496 22752 6560
rect 22816 6496 22832 6560
rect 22896 6496 22912 6560
rect 22976 6496 22992 6560
rect 23056 6496 23064 6560
rect 22744 6046 23064 6496
rect 22744 5810 22786 6046
rect 23022 5810 23064 6046
rect 22744 5472 23064 5810
rect 22744 5408 22752 5472
rect 22816 5408 22832 5472
rect 22896 5408 22912 5472
rect 22976 5408 22992 5472
rect 23056 5408 23064 5472
rect 22744 4384 23064 5408
rect 22744 4320 22752 4384
rect 22816 4320 22832 4384
rect 22896 4320 22912 4384
rect 22976 4320 22992 4384
rect 23056 4320 23064 4384
rect 22744 3296 23064 4320
rect 22744 3232 22752 3296
rect 22816 3232 22832 3296
rect 22896 3232 22912 3296
rect 22976 3232 22992 3296
rect 23056 3232 23064 3296
rect 22744 3046 23064 3232
rect 22744 2810 22786 3046
rect 23022 2810 23064 3046
rect 22744 2208 23064 2810
rect 22744 2144 22752 2208
rect 22816 2144 22832 2208
rect 22896 2144 22912 2208
rect 22976 2144 22992 2208
rect 23056 2144 23064 2208
rect 22744 2128 23064 2144
rect 24244 28864 24564 29424
rect 24244 28800 24252 28864
rect 24316 28800 24332 28864
rect 24396 28800 24412 28864
rect 24476 28800 24492 28864
rect 24556 28800 24564 28864
rect 24244 28546 24564 28800
rect 24244 28310 24286 28546
rect 24522 28310 24564 28546
rect 24244 27776 24564 28310
rect 24244 27712 24252 27776
rect 24316 27712 24332 27776
rect 24396 27712 24412 27776
rect 24476 27712 24492 27776
rect 24556 27712 24564 27776
rect 24244 26688 24564 27712
rect 24244 26624 24252 26688
rect 24316 26624 24332 26688
rect 24396 26624 24412 26688
rect 24476 26624 24492 26688
rect 24556 26624 24564 26688
rect 24244 25600 24564 26624
rect 24244 25536 24252 25600
rect 24316 25546 24332 25600
rect 24396 25546 24412 25600
rect 24476 25546 24492 25600
rect 24556 25536 24564 25600
rect 24244 25310 24286 25536
rect 24522 25310 24564 25536
rect 24244 24512 24564 25310
rect 24244 24448 24252 24512
rect 24316 24448 24332 24512
rect 24396 24448 24412 24512
rect 24476 24448 24492 24512
rect 24556 24448 24564 24512
rect 24244 23424 24564 24448
rect 24244 23360 24252 23424
rect 24316 23360 24332 23424
rect 24396 23360 24412 23424
rect 24476 23360 24492 23424
rect 24556 23360 24564 23424
rect 24244 22546 24564 23360
rect 24244 22336 24286 22546
rect 24522 22336 24564 22546
rect 24244 22272 24252 22336
rect 24316 22272 24332 22310
rect 24396 22272 24412 22310
rect 24476 22272 24492 22310
rect 24556 22272 24564 22336
rect 24244 21248 24564 22272
rect 24244 21184 24252 21248
rect 24316 21184 24332 21248
rect 24396 21184 24412 21248
rect 24476 21184 24492 21248
rect 24556 21184 24564 21248
rect 24244 20160 24564 21184
rect 24244 20096 24252 20160
rect 24316 20096 24332 20160
rect 24396 20096 24412 20160
rect 24476 20096 24492 20160
rect 24556 20096 24564 20160
rect 24244 19546 24564 20096
rect 24244 19310 24286 19546
rect 24522 19310 24564 19546
rect 24244 19072 24564 19310
rect 24244 19008 24252 19072
rect 24316 19008 24332 19072
rect 24396 19008 24412 19072
rect 24476 19008 24492 19072
rect 24556 19008 24564 19072
rect 24244 17984 24564 19008
rect 24244 17920 24252 17984
rect 24316 17920 24332 17984
rect 24396 17920 24412 17984
rect 24476 17920 24492 17984
rect 24556 17920 24564 17984
rect 24244 16896 24564 17920
rect 24244 16832 24252 16896
rect 24316 16832 24332 16896
rect 24396 16832 24412 16896
rect 24476 16832 24492 16896
rect 24556 16832 24564 16896
rect 24244 16546 24564 16832
rect 24244 16310 24286 16546
rect 24522 16310 24564 16546
rect 24244 15808 24564 16310
rect 24244 15744 24252 15808
rect 24316 15744 24332 15808
rect 24396 15744 24412 15808
rect 24476 15744 24492 15808
rect 24556 15744 24564 15808
rect 24244 14720 24564 15744
rect 24244 14656 24252 14720
rect 24316 14656 24332 14720
rect 24396 14656 24412 14720
rect 24476 14656 24492 14720
rect 24556 14656 24564 14720
rect 24244 13632 24564 14656
rect 24244 13568 24252 13632
rect 24316 13568 24332 13632
rect 24396 13568 24412 13632
rect 24476 13568 24492 13632
rect 24556 13568 24564 13632
rect 24244 13546 24564 13568
rect 24244 13310 24286 13546
rect 24522 13310 24564 13546
rect 24244 12544 24564 13310
rect 24244 12480 24252 12544
rect 24316 12480 24332 12544
rect 24396 12480 24412 12544
rect 24476 12480 24492 12544
rect 24556 12480 24564 12544
rect 24244 11456 24564 12480
rect 24244 11392 24252 11456
rect 24316 11392 24332 11456
rect 24396 11392 24412 11456
rect 24476 11392 24492 11456
rect 24556 11392 24564 11456
rect 24244 10546 24564 11392
rect 24244 10368 24286 10546
rect 24522 10368 24564 10546
rect 24244 10304 24252 10368
rect 24316 10304 24332 10310
rect 24396 10304 24412 10310
rect 24476 10304 24492 10310
rect 24556 10304 24564 10368
rect 24244 9280 24564 10304
rect 24244 9216 24252 9280
rect 24316 9216 24332 9280
rect 24396 9216 24412 9280
rect 24476 9216 24492 9280
rect 24556 9216 24564 9280
rect 24244 8192 24564 9216
rect 24244 8128 24252 8192
rect 24316 8128 24332 8192
rect 24396 8128 24412 8192
rect 24476 8128 24492 8192
rect 24556 8128 24564 8192
rect 24244 7546 24564 8128
rect 24244 7310 24286 7546
rect 24522 7310 24564 7546
rect 24244 7104 24564 7310
rect 24244 7040 24252 7104
rect 24316 7040 24332 7104
rect 24396 7040 24412 7104
rect 24476 7040 24492 7104
rect 24556 7040 24564 7104
rect 24244 6016 24564 7040
rect 24244 5952 24252 6016
rect 24316 5952 24332 6016
rect 24396 5952 24412 6016
rect 24476 5952 24492 6016
rect 24556 5952 24564 6016
rect 24244 4928 24564 5952
rect 24244 4864 24252 4928
rect 24316 4864 24332 4928
rect 24396 4864 24412 4928
rect 24476 4864 24492 4928
rect 24556 4864 24564 4928
rect 24244 4546 24564 4864
rect 24244 4310 24286 4546
rect 24522 4310 24564 4546
rect 24244 3840 24564 4310
rect 24244 3776 24252 3840
rect 24316 3776 24332 3840
rect 24396 3776 24412 3840
rect 24476 3776 24492 3840
rect 24556 3776 24564 3840
rect 24244 2752 24564 3776
rect 24244 2688 24252 2752
rect 24316 2688 24332 2752
rect 24396 2688 24412 2752
rect 24476 2688 24492 2752
rect 24556 2688 24564 2752
rect 24244 2128 24564 2688
rect 25744 29408 26064 29424
rect 25744 29344 25752 29408
rect 25816 29344 25832 29408
rect 25896 29344 25912 29408
rect 25976 29344 25992 29408
rect 26056 29344 26064 29408
rect 25744 28320 26064 29344
rect 25744 28256 25752 28320
rect 25816 28256 25832 28320
rect 25896 28256 25912 28320
rect 25976 28256 25992 28320
rect 26056 28256 26064 28320
rect 25744 27232 26064 28256
rect 25744 27168 25752 27232
rect 25816 27168 25832 27232
rect 25896 27168 25912 27232
rect 25976 27168 25992 27232
rect 26056 27168 26064 27232
rect 25744 27046 26064 27168
rect 25744 26810 25786 27046
rect 26022 26810 26064 27046
rect 25744 26144 26064 26810
rect 25744 26080 25752 26144
rect 25816 26080 25832 26144
rect 25896 26080 25912 26144
rect 25976 26080 25992 26144
rect 26056 26080 26064 26144
rect 25744 25056 26064 26080
rect 25744 24992 25752 25056
rect 25816 24992 25832 25056
rect 25896 24992 25912 25056
rect 25976 24992 25992 25056
rect 26056 24992 26064 25056
rect 25744 24046 26064 24992
rect 25744 23968 25786 24046
rect 26022 23968 26064 24046
rect 25744 23904 25752 23968
rect 26056 23904 26064 23968
rect 25744 23810 25786 23904
rect 26022 23810 26064 23904
rect 25744 22880 26064 23810
rect 25744 22816 25752 22880
rect 25816 22816 25832 22880
rect 25896 22816 25912 22880
rect 25976 22816 25992 22880
rect 26056 22816 26064 22880
rect 25744 21792 26064 22816
rect 25744 21728 25752 21792
rect 25816 21728 25832 21792
rect 25896 21728 25912 21792
rect 25976 21728 25992 21792
rect 26056 21728 26064 21792
rect 25744 21046 26064 21728
rect 25744 20810 25786 21046
rect 26022 20810 26064 21046
rect 25744 20704 26064 20810
rect 25744 20640 25752 20704
rect 25816 20640 25832 20704
rect 25896 20640 25912 20704
rect 25976 20640 25992 20704
rect 26056 20640 26064 20704
rect 25744 19616 26064 20640
rect 25744 19552 25752 19616
rect 25816 19552 25832 19616
rect 25896 19552 25912 19616
rect 25976 19552 25992 19616
rect 26056 19552 26064 19616
rect 25744 18528 26064 19552
rect 25744 18464 25752 18528
rect 25816 18464 25832 18528
rect 25896 18464 25912 18528
rect 25976 18464 25992 18528
rect 26056 18464 26064 18528
rect 25744 18046 26064 18464
rect 25744 17810 25786 18046
rect 26022 17810 26064 18046
rect 25744 17440 26064 17810
rect 25744 17376 25752 17440
rect 25816 17376 25832 17440
rect 25896 17376 25912 17440
rect 25976 17376 25992 17440
rect 26056 17376 26064 17440
rect 25744 16352 26064 17376
rect 25744 16288 25752 16352
rect 25816 16288 25832 16352
rect 25896 16288 25912 16352
rect 25976 16288 25992 16352
rect 26056 16288 26064 16352
rect 25744 15264 26064 16288
rect 25744 15200 25752 15264
rect 25816 15200 25832 15264
rect 25896 15200 25912 15264
rect 25976 15200 25992 15264
rect 26056 15200 26064 15264
rect 25744 15046 26064 15200
rect 25744 14810 25786 15046
rect 26022 14810 26064 15046
rect 25744 14176 26064 14810
rect 25744 14112 25752 14176
rect 25816 14112 25832 14176
rect 25896 14112 25912 14176
rect 25976 14112 25992 14176
rect 26056 14112 26064 14176
rect 25744 13088 26064 14112
rect 25744 13024 25752 13088
rect 25816 13024 25832 13088
rect 25896 13024 25912 13088
rect 25976 13024 25992 13088
rect 26056 13024 26064 13088
rect 25744 12046 26064 13024
rect 25744 12000 25786 12046
rect 26022 12000 26064 12046
rect 25744 11936 25752 12000
rect 26056 11936 26064 12000
rect 25744 11810 25786 11936
rect 26022 11810 26064 11936
rect 25744 10912 26064 11810
rect 25744 10848 25752 10912
rect 25816 10848 25832 10912
rect 25896 10848 25912 10912
rect 25976 10848 25992 10912
rect 26056 10848 26064 10912
rect 25744 9824 26064 10848
rect 25744 9760 25752 9824
rect 25816 9760 25832 9824
rect 25896 9760 25912 9824
rect 25976 9760 25992 9824
rect 26056 9760 26064 9824
rect 25744 9046 26064 9760
rect 25744 8810 25786 9046
rect 26022 8810 26064 9046
rect 25744 8736 26064 8810
rect 25744 8672 25752 8736
rect 25816 8672 25832 8736
rect 25896 8672 25912 8736
rect 25976 8672 25992 8736
rect 26056 8672 26064 8736
rect 25744 7648 26064 8672
rect 25744 7584 25752 7648
rect 25816 7584 25832 7648
rect 25896 7584 25912 7648
rect 25976 7584 25992 7648
rect 26056 7584 26064 7648
rect 25744 6560 26064 7584
rect 25744 6496 25752 6560
rect 25816 6496 25832 6560
rect 25896 6496 25912 6560
rect 25976 6496 25992 6560
rect 26056 6496 26064 6560
rect 25744 6046 26064 6496
rect 25744 5810 25786 6046
rect 26022 5810 26064 6046
rect 25744 5472 26064 5810
rect 25744 5408 25752 5472
rect 25816 5408 25832 5472
rect 25896 5408 25912 5472
rect 25976 5408 25992 5472
rect 26056 5408 26064 5472
rect 25744 4384 26064 5408
rect 25744 4320 25752 4384
rect 25816 4320 25832 4384
rect 25896 4320 25912 4384
rect 25976 4320 25992 4384
rect 26056 4320 26064 4384
rect 25744 3296 26064 4320
rect 25744 3232 25752 3296
rect 25816 3232 25832 3296
rect 25896 3232 25912 3296
rect 25976 3232 25992 3296
rect 26056 3232 26064 3296
rect 25744 3046 26064 3232
rect 25744 2810 25786 3046
rect 26022 2810 26064 3046
rect 25744 2208 26064 2810
rect 25744 2144 25752 2208
rect 25816 2144 25832 2208
rect 25896 2144 25912 2208
rect 25976 2144 25992 2208
rect 26056 2144 26064 2208
rect 25744 2128 26064 2144
rect 27244 28864 27564 29424
rect 27244 28800 27252 28864
rect 27316 28800 27332 28864
rect 27396 28800 27412 28864
rect 27476 28800 27492 28864
rect 27556 28800 27564 28864
rect 27244 28546 27564 28800
rect 27244 28310 27286 28546
rect 27522 28310 27564 28546
rect 27244 27776 27564 28310
rect 27244 27712 27252 27776
rect 27316 27712 27332 27776
rect 27396 27712 27412 27776
rect 27476 27712 27492 27776
rect 27556 27712 27564 27776
rect 27244 26688 27564 27712
rect 27244 26624 27252 26688
rect 27316 26624 27332 26688
rect 27396 26624 27412 26688
rect 27476 26624 27492 26688
rect 27556 26624 27564 26688
rect 27244 25600 27564 26624
rect 27244 25536 27252 25600
rect 27316 25546 27332 25600
rect 27396 25546 27412 25600
rect 27476 25546 27492 25600
rect 27556 25536 27564 25600
rect 27244 25310 27286 25536
rect 27522 25310 27564 25536
rect 27244 24512 27564 25310
rect 27244 24448 27252 24512
rect 27316 24448 27332 24512
rect 27396 24448 27412 24512
rect 27476 24448 27492 24512
rect 27556 24448 27564 24512
rect 27244 23424 27564 24448
rect 27244 23360 27252 23424
rect 27316 23360 27332 23424
rect 27396 23360 27412 23424
rect 27476 23360 27492 23424
rect 27556 23360 27564 23424
rect 27244 22546 27564 23360
rect 27244 22336 27286 22546
rect 27522 22336 27564 22546
rect 27244 22272 27252 22336
rect 27316 22272 27332 22310
rect 27396 22272 27412 22310
rect 27476 22272 27492 22310
rect 27556 22272 27564 22336
rect 27244 21248 27564 22272
rect 27244 21184 27252 21248
rect 27316 21184 27332 21248
rect 27396 21184 27412 21248
rect 27476 21184 27492 21248
rect 27556 21184 27564 21248
rect 27244 20160 27564 21184
rect 27244 20096 27252 20160
rect 27316 20096 27332 20160
rect 27396 20096 27412 20160
rect 27476 20096 27492 20160
rect 27556 20096 27564 20160
rect 27244 19546 27564 20096
rect 27244 19310 27286 19546
rect 27522 19310 27564 19546
rect 27244 19072 27564 19310
rect 27244 19008 27252 19072
rect 27316 19008 27332 19072
rect 27396 19008 27412 19072
rect 27476 19008 27492 19072
rect 27556 19008 27564 19072
rect 27244 17984 27564 19008
rect 27244 17920 27252 17984
rect 27316 17920 27332 17984
rect 27396 17920 27412 17984
rect 27476 17920 27492 17984
rect 27556 17920 27564 17984
rect 27244 16896 27564 17920
rect 27244 16832 27252 16896
rect 27316 16832 27332 16896
rect 27396 16832 27412 16896
rect 27476 16832 27492 16896
rect 27556 16832 27564 16896
rect 27244 16546 27564 16832
rect 27244 16310 27286 16546
rect 27522 16310 27564 16546
rect 27244 15808 27564 16310
rect 27244 15744 27252 15808
rect 27316 15744 27332 15808
rect 27396 15744 27412 15808
rect 27476 15744 27492 15808
rect 27556 15744 27564 15808
rect 27244 14720 27564 15744
rect 27244 14656 27252 14720
rect 27316 14656 27332 14720
rect 27396 14656 27412 14720
rect 27476 14656 27492 14720
rect 27556 14656 27564 14720
rect 27244 13632 27564 14656
rect 27244 13568 27252 13632
rect 27316 13568 27332 13632
rect 27396 13568 27412 13632
rect 27476 13568 27492 13632
rect 27556 13568 27564 13632
rect 27244 13546 27564 13568
rect 27244 13310 27286 13546
rect 27522 13310 27564 13546
rect 27244 12544 27564 13310
rect 27244 12480 27252 12544
rect 27316 12480 27332 12544
rect 27396 12480 27412 12544
rect 27476 12480 27492 12544
rect 27556 12480 27564 12544
rect 27244 11456 27564 12480
rect 27244 11392 27252 11456
rect 27316 11392 27332 11456
rect 27396 11392 27412 11456
rect 27476 11392 27492 11456
rect 27556 11392 27564 11456
rect 27244 10546 27564 11392
rect 27244 10368 27286 10546
rect 27522 10368 27564 10546
rect 27244 10304 27252 10368
rect 27316 10304 27332 10310
rect 27396 10304 27412 10310
rect 27476 10304 27492 10310
rect 27556 10304 27564 10368
rect 27244 9280 27564 10304
rect 27244 9216 27252 9280
rect 27316 9216 27332 9280
rect 27396 9216 27412 9280
rect 27476 9216 27492 9280
rect 27556 9216 27564 9280
rect 27244 8192 27564 9216
rect 27244 8128 27252 8192
rect 27316 8128 27332 8192
rect 27396 8128 27412 8192
rect 27476 8128 27492 8192
rect 27556 8128 27564 8192
rect 27244 7546 27564 8128
rect 27244 7310 27286 7546
rect 27522 7310 27564 7546
rect 27244 7104 27564 7310
rect 27244 7040 27252 7104
rect 27316 7040 27332 7104
rect 27396 7040 27412 7104
rect 27476 7040 27492 7104
rect 27556 7040 27564 7104
rect 27244 6016 27564 7040
rect 27244 5952 27252 6016
rect 27316 5952 27332 6016
rect 27396 5952 27412 6016
rect 27476 5952 27492 6016
rect 27556 5952 27564 6016
rect 27244 4928 27564 5952
rect 27244 4864 27252 4928
rect 27316 4864 27332 4928
rect 27396 4864 27412 4928
rect 27476 4864 27492 4928
rect 27556 4864 27564 4928
rect 27244 4546 27564 4864
rect 27244 4310 27286 4546
rect 27522 4310 27564 4546
rect 27244 3840 27564 4310
rect 27244 3776 27252 3840
rect 27316 3776 27332 3840
rect 27396 3776 27412 3840
rect 27476 3776 27492 3840
rect 27556 3776 27564 3840
rect 27244 2752 27564 3776
rect 27244 2688 27252 2752
rect 27316 2688 27332 2752
rect 27396 2688 27412 2752
rect 27476 2688 27492 2752
rect 27556 2688 27564 2752
rect 27244 2128 27564 2688
<< via4 >>
rect 1786 26810 2022 27046
rect 1786 23968 2022 24046
rect 1786 23904 1816 23968
rect 1816 23904 1832 23968
rect 1832 23904 1896 23968
rect 1896 23904 1912 23968
rect 1912 23904 1976 23968
rect 1976 23904 1992 23968
rect 1992 23904 2022 23968
rect 1786 23810 2022 23904
rect 1786 20810 2022 21046
rect 1786 17810 2022 18046
rect 1786 14810 2022 15046
rect 1786 12000 2022 12046
rect 1786 11936 1816 12000
rect 1816 11936 1832 12000
rect 1832 11936 1896 12000
rect 1896 11936 1912 12000
rect 1912 11936 1976 12000
rect 1976 11936 1992 12000
rect 1992 11936 2022 12000
rect 1786 11810 2022 11936
rect 1786 8810 2022 9046
rect 1786 5810 2022 6046
rect 1786 2810 2022 3046
rect 3286 28310 3522 28546
rect 3286 25536 3316 25546
rect 3316 25536 3332 25546
rect 3332 25536 3396 25546
rect 3396 25536 3412 25546
rect 3412 25536 3476 25546
rect 3476 25536 3492 25546
rect 3492 25536 3522 25546
rect 3286 25310 3522 25536
rect 3286 22336 3522 22546
rect 3286 22310 3316 22336
rect 3316 22310 3332 22336
rect 3332 22310 3396 22336
rect 3396 22310 3412 22336
rect 3412 22310 3476 22336
rect 3476 22310 3492 22336
rect 3492 22310 3522 22336
rect 3286 19310 3522 19546
rect 3286 16310 3522 16546
rect 3286 13310 3522 13546
rect 3286 10368 3522 10546
rect 3286 10310 3316 10368
rect 3316 10310 3332 10368
rect 3332 10310 3396 10368
rect 3396 10310 3412 10368
rect 3412 10310 3476 10368
rect 3476 10310 3492 10368
rect 3492 10310 3522 10368
rect 3286 7310 3522 7546
rect 3286 4310 3522 4546
rect 4786 26810 5022 27046
rect 4786 23968 5022 24046
rect 4786 23904 4816 23968
rect 4816 23904 4832 23968
rect 4832 23904 4896 23968
rect 4896 23904 4912 23968
rect 4912 23904 4976 23968
rect 4976 23904 4992 23968
rect 4992 23904 5022 23968
rect 4786 23810 5022 23904
rect 4786 20810 5022 21046
rect 4786 17810 5022 18046
rect 4786 14810 5022 15046
rect 4786 12000 5022 12046
rect 4786 11936 4816 12000
rect 4816 11936 4832 12000
rect 4832 11936 4896 12000
rect 4896 11936 4912 12000
rect 4912 11936 4976 12000
rect 4976 11936 4992 12000
rect 4992 11936 5022 12000
rect 4786 11810 5022 11936
rect 4786 8810 5022 9046
rect 4786 5810 5022 6046
rect 4786 2810 5022 3046
rect 6286 28310 6522 28546
rect 6286 25536 6316 25546
rect 6316 25536 6332 25546
rect 6332 25536 6396 25546
rect 6396 25536 6412 25546
rect 6412 25536 6476 25546
rect 6476 25536 6492 25546
rect 6492 25536 6522 25546
rect 6286 25310 6522 25536
rect 6286 22336 6522 22546
rect 6286 22310 6316 22336
rect 6316 22310 6332 22336
rect 6332 22310 6396 22336
rect 6396 22310 6412 22336
rect 6412 22310 6476 22336
rect 6476 22310 6492 22336
rect 6492 22310 6522 22336
rect 6286 19310 6522 19546
rect 6286 16310 6522 16546
rect 6286 13310 6522 13546
rect 6286 10368 6522 10546
rect 6286 10310 6316 10368
rect 6316 10310 6332 10368
rect 6332 10310 6396 10368
rect 6396 10310 6412 10368
rect 6412 10310 6476 10368
rect 6476 10310 6492 10368
rect 6492 10310 6522 10368
rect 6286 7310 6522 7546
rect 6286 4310 6522 4546
rect 7786 26810 8022 27046
rect 7786 23968 8022 24046
rect 7786 23904 7816 23968
rect 7816 23904 7832 23968
rect 7832 23904 7896 23968
rect 7896 23904 7912 23968
rect 7912 23904 7976 23968
rect 7976 23904 7992 23968
rect 7992 23904 8022 23968
rect 7786 23810 8022 23904
rect 7786 20810 8022 21046
rect 7786 17810 8022 18046
rect 7786 14810 8022 15046
rect 7786 12000 8022 12046
rect 7786 11936 7816 12000
rect 7816 11936 7832 12000
rect 7832 11936 7896 12000
rect 7896 11936 7912 12000
rect 7912 11936 7976 12000
rect 7976 11936 7992 12000
rect 7992 11936 8022 12000
rect 7786 11810 8022 11936
rect 7786 8810 8022 9046
rect 7786 5810 8022 6046
rect 7786 2810 8022 3046
rect 9286 28310 9522 28546
rect 9286 25536 9316 25546
rect 9316 25536 9332 25546
rect 9332 25536 9396 25546
rect 9396 25536 9412 25546
rect 9412 25536 9476 25546
rect 9476 25536 9492 25546
rect 9492 25536 9522 25546
rect 9286 25310 9522 25536
rect 9286 22336 9522 22546
rect 9286 22310 9316 22336
rect 9316 22310 9332 22336
rect 9332 22310 9396 22336
rect 9396 22310 9412 22336
rect 9412 22310 9476 22336
rect 9476 22310 9492 22336
rect 9492 22310 9522 22336
rect 9286 19310 9522 19546
rect 9286 16310 9522 16546
rect 9286 13310 9522 13546
rect 9286 10368 9522 10546
rect 9286 10310 9316 10368
rect 9316 10310 9332 10368
rect 9332 10310 9396 10368
rect 9396 10310 9412 10368
rect 9412 10310 9476 10368
rect 9476 10310 9492 10368
rect 9492 10310 9522 10368
rect 9286 7310 9522 7546
rect 9286 4310 9522 4546
rect 10786 26810 11022 27046
rect 10786 23968 11022 24046
rect 10786 23904 10816 23968
rect 10816 23904 10832 23968
rect 10832 23904 10896 23968
rect 10896 23904 10912 23968
rect 10912 23904 10976 23968
rect 10976 23904 10992 23968
rect 10992 23904 11022 23968
rect 10786 23810 11022 23904
rect 10786 20810 11022 21046
rect 10786 17810 11022 18046
rect 10786 14810 11022 15046
rect 10786 12000 11022 12046
rect 10786 11936 10816 12000
rect 10816 11936 10832 12000
rect 10832 11936 10896 12000
rect 10896 11936 10912 12000
rect 10912 11936 10976 12000
rect 10976 11936 10992 12000
rect 10992 11936 11022 12000
rect 10786 11810 11022 11936
rect 10786 8810 11022 9046
rect 10786 5810 11022 6046
rect 10786 2810 11022 3046
rect 12286 28310 12522 28546
rect 12286 25536 12316 25546
rect 12316 25536 12332 25546
rect 12332 25536 12396 25546
rect 12396 25536 12412 25546
rect 12412 25536 12476 25546
rect 12476 25536 12492 25546
rect 12492 25536 12522 25546
rect 12286 25310 12522 25536
rect 12286 22336 12522 22546
rect 12286 22310 12316 22336
rect 12316 22310 12332 22336
rect 12332 22310 12396 22336
rect 12396 22310 12412 22336
rect 12412 22310 12476 22336
rect 12476 22310 12492 22336
rect 12492 22310 12522 22336
rect 12286 19310 12522 19546
rect 12286 16310 12522 16546
rect 12286 13310 12522 13546
rect 12286 10368 12522 10546
rect 12286 10310 12316 10368
rect 12316 10310 12332 10368
rect 12332 10310 12396 10368
rect 12396 10310 12412 10368
rect 12412 10310 12476 10368
rect 12476 10310 12492 10368
rect 12492 10310 12522 10368
rect 12286 7310 12522 7546
rect 12286 4310 12522 4546
rect 13786 26810 14022 27046
rect 13786 23968 14022 24046
rect 13786 23904 13816 23968
rect 13816 23904 13832 23968
rect 13832 23904 13896 23968
rect 13896 23904 13912 23968
rect 13912 23904 13976 23968
rect 13976 23904 13992 23968
rect 13992 23904 14022 23968
rect 13786 23810 14022 23904
rect 13786 20810 14022 21046
rect 13786 17810 14022 18046
rect 13786 14810 14022 15046
rect 13786 12000 14022 12046
rect 13786 11936 13816 12000
rect 13816 11936 13832 12000
rect 13832 11936 13896 12000
rect 13896 11936 13912 12000
rect 13912 11936 13976 12000
rect 13976 11936 13992 12000
rect 13992 11936 14022 12000
rect 13786 11810 14022 11936
rect 13786 8810 14022 9046
rect 13786 5810 14022 6046
rect 13786 2810 14022 3046
rect 15286 28310 15522 28546
rect 15286 25536 15316 25546
rect 15316 25536 15332 25546
rect 15332 25536 15396 25546
rect 15396 25536 15412 25546
rect 15412 25536 15476 25546
rect 15476 25536 15492 25546
rect 15492 25536 15522 25546
rect 15286 25310 15522 25536
rect 15286 22336 15522 22546
rect 15286 22310 15316 22336
rect 15316 22310 15332 22336
rect 15332 22310 15396 22336
rect 15396 22310 15412 22336
rect 15412 22310 15476 22336
rect 15476 22310 15492 22336
rect 15492 22310 15522 22336
rect 15286 19310 15522 19546
rect 15286 16310 15522 16546
rect 15286 13310 15522 13546
rect 15286 10368 15522 10546
rect 15286 10310 15316 10368
rect 15316 10310 15332 10368
rect 15332 10310 15396 10368
rect 15396 10310 15412 10368
rect 15412 10310 15476 10368
rect 15476 10310 15492 10368
rect 15492 10310 15522 10368
rect 15286 7310 15522 7546
rect 15286 4310 15522 4546
rect 16786 26810 17022 27046
rect 16786 23968 17022 24046
rect 16786 23904 16816 23968
rect 16816 23904 16832 23968
rect 16832 23904 16896 23968
rect 16896 23904 16912 23968
rect 16912 23904 16976 23968
rect 16976 23904 16992 23968
rect 16992 23904 17022 23968
rect 16786 23810 17022 23904
rect 16786 20810 17022 21046
rect 16786 17810 17022 18046
rect 16786 14810 17022 15046
rect 16786 12000 17022 12046
rect 16786 11936 16816 12000
rect 16816 11936 16832 12000
rect 16832 11936 16896 12000
rect 16896 11936 16912 12000
rect 16912 11936 16976 12000
rect 16976 11936 16992 12000
rect 16992 11936 17022 12000
rect 16786 11810 17022 11936
rect 16786 8810 17022 9046
rect 16786 5810 17022 6046
rect 16786 2810 17022 3046
rect 18286 28310 18522 28546
rect 18286 25536 18316 25546
rect 18316 25536 18332 25546
rect 18332 25536 18396 25546
rect 18396 25536 18412 25546
rect 18412 25536 18476 25546
rect 18476 25536 18492 25546
rect 18492 25536 18522 25546
rect 18286 25310 18522 25536
rect 18286 22336 18522 22546
rect 18286 22310 18316 22336
rect 18316 22310 18332 22336
rect 18332 22310 18396 22336
rect 18396 22310 18412 22336
rect 18412 22310 18476 22336
rect 18476 22310 18492 22336
rect 18492 22310 18522 22336
rect 18286 19310 18522 19546
rect 18286 16310 18522 16546
rect 19786 26810 20022 27046
rect 19786 23968 20022 24046
rect 19786 23904 19816 23968
rect 19816 23904 19832 23968
rect 19832 23904 19896 23968
rect 19896 23904 19912 23968
rect 19912 23904 19976 23968
rect 19976 23904 19992 23968
rect 19992 23904 20022 23968
rect 19786 23810 20022 23904
rect 19786 20810 20022 21046
rect 19786 17810 20022 18046
rect 19786 14810 20022 15046
rect 18286 13310 18522 13546
rect 18286 10368 18522 10546
rect 18286 10310 18316 10368
rect 18316 10310 18332 10368
rect 18332 10310 18396 10368
rect 18396 10310 18412 10368
rect 18412 10310 18476 10368
rect 18476 10310 18492 10368
rect 18492 10310 18522 10368
rect 19786 12000 20022 12046
rect 19786 11936 19816 12000
rect 19816 11936 19832 12000
rect 19832 11936 19896 12000
rect 19896 11936 19912 12000
rect 19912 11936 19976 12000
rect 19976 11936 19992 12000
rect 19992 11936 20022 12000
rect 19786 11810 20022 11936
rect 18286 7310 18522 7546
rect 18286 4310 18522 4546
rect 19786 8810 20022 9046
rect 19786 5810 20022 6046
rect 19786 2810 20022 3046
rect 21286 28310 21522 28546
rect 21286 25536 21316 25546
rect 21316 25536 21332 25546
rect 21332 25536 21396 25546
rect 21396 25536 21412 25546
rect 21412 25536 21476 25546
rect 21476 25536 21492 25546
rect 21492 25536 21522 25546
rect 21286 25310 21522 25536
rect 21286 22336 21522 22546
rect 21286 22310 21316 22336
rect 21316 22310 21332 22336
rect 21332 22310 21396 22336
rect 21396 22310 21412 22336
rect 21412 22310 21476 22336
rect 21476 22310 21492 22336
rect 21492 22310 21522 22336
rect 21286 19310 21522 19546
rect 21286 16310 21522 16546
rect 21286 13310 21522 13546
rect 21286 10368 21522 10546
rect 21286 10310 21316 10368
rect 21316 10310 21332 10368
rect 21332 10310 21396 10368
rect 21396 10310 21412 10368
rect 21412 10310 21476 10368
rect 21476 10310 21492 10368
rect 21492 10310 21522 10368
rect 21286 7310 21522 7546
rect 21286 4310 21522 4546
rect 22786 26810 23022 27046
rect 22786 23968 23022 24046
rect 22786 23904 22816 23968
rect 22816 23904 22832 23968
rect 22832 23904 22896 23968
rect 22896 23904 22912 23968
rect 22912 23904 22976 23968
rect 22976 23904 22992 23968
rect 22992 23904 23022 23968
rect 22786 23810 23022 23904
rect 22786 20810 23022 21046
rect 22786 17810 23022 18046
rect 22786 14810 23022 15046
rect 22786 12000 23022 12046
rect 22786 11936 22816 12000
rect 22816 11936 22832 12000
rect 22832 11936 22896 12000
rect 22896 11936 22912 12000
rect 22912 11936 22976 12000
rect 22976 11936 22992 12000
rect 22992 11936 23022 12000
rect 22786 11810 23022 11936
rect 22786 8810 23022 9046
rect 22786 5810 23022 6046
rect 22786 2810 23022 3046
rect 24286 28310 24522 28546
rect 24286 25536 24316 25546
rect 24316 25536 24332 25546
rect 24332 25536 24396 25546
rect 24396 25536 24412 25546
rect 24412 25536 24476 25546
rect 24476 25536 24492 25546
rect 24492 25536 24522 25546
rect 24286 25310 24522 25536
rect 24286 22336 24522 22546
rect 24286 22310 24316 22336
rect 24316 22310 24332 22336
rect 24332 22310 24396 22336
rect 24396 22310 24412 22336
rect 24412 22310 24476 22336
rect 24476 22310 24492 22336
rect 24492 22310 24522 22336
rect 24286 19310 24522 19546
rect 24286 16310 24522 16546
rect 24286 13310 24522 13546
rect 24286 10368 24522 10546
rect 24286 10310 24316 10368
rect 24316 10310 24332 10368
rect 24332 10310 24396 10368
rect 24396 10310 24412 10368
rect 24412 10310 24476 10368
rect 24476 10310 24492 10368
rect 24492 10310 24522 10368
rect 24286 7310 24522 7546
rect 24286 4310 24522 4546
rect 25786 26810 26022 27046
rect 25786 23968 26022 24046
rect 25786 23904 25816 23968
rect 25816 23904 25832 23968
rect 25832 23904 25896 23968
rect 25896 23904 25912 23968
rect 25912 23904 25976 23968
rect 25976 23904 25992 23968
rect 25992 23904 26022 23968
rect 25786 23810 26022 23904
rect 25786 20810 26022 21046
rect 25786 17810 26022 18046
rect 25786 14810 26022 15046
rect 25786 12000 26022 12046
rect 25786 11936 25816 12000
rect 25816 11936 25832 12000
rect 25832 11936 25896 12000
rect 25896 11936 25912 12000
rect 25912 11936 25976 12000
rect 25976 11936 25992 12000
rect 25992 11936 26022 12000
rect 25786 11810 26022 11936
rect 25786 8810 26022 9046
rect 25786 5810 26022 6046
rect 25786 2810 26022 3046
rect 27286 28310 27522 28546
rect 27286 25536 27316 25546
rect 27316 25536 27332 25546
rect 27332 25536 27396 25546
rect 27396 25536 27412 25546
rect 27412 25536 27476 25546
rect 27476 25536 27492 25546
rect 27492 25536 27522 25546
rect 27286 25310 27522 25536
rect 27286 22336 27522 22546
rect 27286 22310 27316 22336
rect 27316 22310 27332 22336
rect 27332 22310 27396 22336
rect 27396 22310 27412 22336
rect 27412 22310 27476 22336
rect 27476 22310 27492 22336
rect 27492 22310 27522 22336
rect 27286 19310 27522 19546
rect 27286 16310 27522 16546
rect 27286 13310 27522 13546
rect 27286 10368 27522 10546
rect 27286 10310 27316 10368
rect 27316 10310 27332 10368
rect 27332 10310 27396 10368
rect 27396 10310 27412 10368
rect 27412 10310 27476 10368
rect 27476 10310 27492 10368
rect 27492 10310 27522 10368
rect 27286 7310 27522 7546
rect 27286 4310 27522 4546
<< metal5 >>
rect 1104 28546 28336 28588
rect 1104 28310 3286 28546
rect 3522 28310 6286 28546
rect 6522 28310 9286 28546
rect 9522 28310 12286 28546
rect 12522 28310 15286 28546
rect 15522 28310 18286 28546
rect 18522 28310 21286 28546
rect 21522 28310 24286 28546
rect 24522 28310 27286 28546
rect 27522 28310 28336 28546
rect 1104 28268 28336 28310
rect 1104 27046 28336 27088
rect 1104 26810 1786 27046
rect 2022 26810 4786 27046
rect 5022 26810 7786 27046
rect 8022 26810 10786 27046
rect 11022 26810 13786 27046
rect 14022 26810 16786 27046
rect 17022 26810 19786 27046
rect 20022 26810 22786 27046
rect 23022 26810 25786 27046
rect 26022 26810 28336 27046
rect 1104 26768 28336 26810
rect 1104 25546 28336 25588
rect 1104 25310 3286 25546
rect 3522 25310 6286 25546
rect 6522 25310 9286 25546
rect 9522 25310 12286 25546
rect 12522 25310 15286 25546
rect 15522 25310 18286 25546
rect 18522 25310 21286 25546
rect 21522 25310 24286 25546
rect 24522 25310 27286 25546
rect 27522 25310 28336 25546
rect 1104 25268 28336 25310
rect 1104 24046 28336 24088
rect 1104 23810 1786 24046
rect 2022 23810 4786 24046
rect 5022 23810 7786 24046
rect 8022 23810 10786 24046
rect 11022 23810 13786 24046
rect 14022 23810 16786 24046
rect 17022 23810 19786 24046
rect 20022 23810 22786 24046
rect 23022 23810 25786 24046
rect 26022 23810 28336 24046
rect 1104 23768 28336 23810
rect 1104 22546 28336 22588
rect 1104 22310 3286 22546
rect 3522 22310 6286 22546
rect 6522 22310 9286 22546
rect 9522 22310 12286 22546
rect 12522 22310 15286 22546
rect 15522 22310 18286 22546
rect 18522 22310 21286 22546
rect 21522 22310 24286 22546
rect 24522 22310 27286 22546
rect 27522 22310 28336 22546
rect 1104 22268 28336 22310
rect 1104 21046 28336 21088
rect 1104 20810 1786 21046
rect 2022 20810 4786 21046
rect 5022 20810 7786 21046
rect 8022 20810 10786 21046
rect 11022 20810 13786 21046
rect 14022 20810 16786 21046
rect 17022 20810 19786 21046
rect 20022 20810 22786 21046
rect 23022 20810 25786 21046
rect 26022 20810 28336 21046
rect 1104 20768 28336 20810
rect 1104 19546 28336 19588
rect 1104 19310 3286 19546
rect 3522 19310 6286 19546
rect 6522 19310 9286 19546
rect 9522 19310 12286 19546
rect 12522 19310 15286 19546
rect 15522 19310 18286 19546
rect 18522 19310 21286 19546
rect 21522 19310 24286 19546
rect 24522 19310 27286 19546
rect 27522 19310 28336 19546
rect 1104 19268 28336 19310
rect 1104 18046 28336 18088
rect 1104 17810 1786 18046
rect 2022 17810 4786 18046
rect 5022 17810 7786 18046
rect 8022 17810 10786 18046
rect 11022 17810 13786 18046
rect 14022 17810 16786 18046
rect 17022 17810 19786 18046
rect 20022 17810 22786 18046
rect 23022 17810 25786 18046
rect 26022 17810 28336 18046
rect 1104 17768 28336 17810
rect 1104 16546 28336 16588
rect 1104 16310 3286 16546
rect 3522 16310 6286 16546
rect 6522 16310 9286 16546
rect 9522 16310 12286 16546
rect 12522 16310 15286 16546
rect 15522 16310 18286 16546
rect 18522 16310 21286 16546
rect 21522 16310 24286 16546
rect 24522 16310 27286 16546
rect 27522 16310 28336 16546
rect 1104 16268 28336 16310
rect 1104 15046 28336 15088
rect 1104 14810 1786 15046
rect 2022 14810 4786 15046
rect 5022 14810 7786 15046
rect 8022 14810 10786 15046
rect 11022 14810 13786 15046
rect 14022 14810 16786 15046
rect 17022 14810 19786 15046
rect 20022 14810 22786 15046
rect 23022 14810 25786 15046
rect 26022 14810 28336 15046
rect 1104 14768 28336 14810
rect 1104 13546 28336 13588
rect 1104 13310 3286 13546
rect 3522 13310 6286 13546
rect 6522 13310 9286 13546
rect 9522 13310 12286 13546
rect 12522 13310 15286 13546
rect 15522 13310 18286 13546
rect 18522 13310 21286 13546
rect 21522 13310 24286 13546
rect 24522 13310 27286 13546
rect 27522 13310 28336 13546
rect 1104 13268 28336 13310
rect 1104 12046 28336 12088
rect 1104 11810 1786 12046
rect 2022 11810 4786 12046
rect 5022 11810 7786 12046
rect 8022 11810 10786 12046
rect 11022 11810 13786 12046
rect 14022 11810 16786 12046
rect 17022 11810 19786 12046
rect 20022 11810 22786 12046
rect 23022 11810 25786 12046
rect 26022 11810 28336 12046
rect 1104 11768 28336 11810
rect 1104 10546 28336 10588
rect 1104 10310 3286 10546
rect 3522 10310 6286 10546
rect 6522 10310 9286 10546
rect 9522 10310 12286 10546
rect 12522 10310 15286 10546
rect 15522 10310 18286 10546
rect 18522 10310 21286 10546
rect 21522 10310 24286 10546
rect 24522 10310 27286 10546
rect 27522 10310 28336 10546
rect 1104 10268 28336 10310
rect 1104 9046 28336 9088
rect 1104 8810 1786 9046
rect 2022 8810 4786 9046
rect 5022 8810 7786 9046
rect 8022 8810 10786 9046
rect 11022 8810 13786 9046
rect 14022 8810 16786 9046
rect 17022 8810 19786 9046
rect 20022 8810 22786 9046
rect 23022 8810 25786 9046
rect 26022 8810 28336 9046
rect 1104 8768 28336 8810
rect 1104 7546 28336 7588
rect 1104 7310 3286 7546
rect 3522 7310 6286 7546
rect 6522 7310 9286 7546
rect 9522 7310 12286 7546
rect 12522 7310 15286 7546
rect 15522 7310 18286 7546
rect 18522 7310 21286 7546
rect 21522 7310 24286 7546
rect 24522 7310 27286 7546
rect 27522 7310 28336 7546
rect 1104 7268 28336 7310
rect 1104 6046 28336 6088
rect 1104 5810 1786 6046
rect 2022 5810 4786 6046
rect 5022 5810 7786 6046
rect 8022 5810 10786 6046
rect 11022 5810 13786 6046
rect 14022 5810 16786 6046
rect 17022 5810 19786 6046
rect 20022 5810 22786 6046
rect 23022 5810 25786 6046
rect 26022 5810 28336 6046
rect 1104 5768 28336 5810
rect 1104 4546 28336 4588
rect 1104 4310 3286 4546
rect 3522 4310 6286 4546
rect 6522 4310 9286 4546
rect 9522 4310 12286 4546
rect 12522 4310 15286 4546
rect 15522 4310 18286 4546
rect 18522 4310 21286 4546
rect 21522 4310 24286 4546
rect 24522 4310 27286 4546
rect 27522 4310 28336 4546
rect 1104 4268 28336 4310
rect 1104 3046 28336 3088
rect 1104 2810 1786 3046
rect 2022 2810 4786 3046
rect 5022 2810 7786 3046
rect 8022 2810 10786 3046
rect 11022 2810 13786 3046
rect 14022 2810 16786 3046
rect 17022 2810 19786 3046
rect 20022 2810 22786 3046
rect 23022 2810 25786 3046
rect 26022 2810 28336 3046
rect 1104 2768 28336 2810
use sky130_fd_sc_hd__decap_12  FILLER_2_15 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1597341371
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1597341371
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1597341371
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1597341371
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1597341371
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1597341371
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1597341371
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1597341371
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1597341371
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1597341371
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1597341371
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1597341371
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1597341371
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1597341371
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1597341371
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1597341371
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1597341371
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_68
timestamp 1597341371
transform 1 0 7360 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1597341371
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1597341371
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63
timestamp 1597341371
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__B home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1597341371
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1597341371
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1597341371
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1597341371
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__B
timestamp 1597341371
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_78
timestamp 1597341371
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1597341371
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1597341371
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1597341371
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_82
timestamp 1597341371
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1597341371
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1597341371
transform 1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A1
timestamp 1597341371
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__B1_N
timestamp 1597341371
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__D
timestamp 1597341371
transform 1 0 8832 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_86
timestamp 1597341371
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1597341371
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1597341371
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1597341371
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1597341371
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1597341371
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A2
timestamp 1597341371
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__RESET_B
timestamp 1597341371
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__CLK
timestamp 1597341371
transform 1 0 9200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1597341371
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1597341371
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1597341371
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1597341371
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _149_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_97 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1597341371
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _290_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10120 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__a21bo_4  _206_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 9568 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1597341371
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1597341371
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1597341371
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__D
timestamp 1597341371
transform 1 0 10396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__CLK
timestamp 1597341371
transform 1 0 10948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _203_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10948 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1597341371
transform 1 0 11868 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1597341371
transform 1 0 11500 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116
timestamp 1597341371
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1597341371
transform 1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__C
timestamp 1597341371
transform 1 0 11316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 1597341371
transform 1 0 12236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1597341371
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1597341371
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1597341371
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__C
timestamp 1597341371
transform 1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1597341371
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1597341371
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1597341371
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_125
timestamp 1597341371
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_128
timestamp 1597341371
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1597341371
transform 1 0 12972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1597341371
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__B1
timestamp 1597341371
transform 1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1597341371
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1597341371
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1597341371
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A2
timestamp 1597341371
transform 1 0 13064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__D
timestamp 1597341371
transform 1 0 13064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1597341371
transform 1 0 13616 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_136
timestamp 1597341371
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__CLK
timestamp 1597341371
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_147
timestamp 1597341371
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_143
timestamp 1597341371
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1597341371
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1597341371
transform 1 0 14812 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A1
timestamp 1597341371
transform 1 0 14444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__RESET_B
timestamp 1597341371
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _195_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 13800 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _289_
timestamp 1597341371
transform 1 0 13708 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__a21oi_4  _202_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 13064 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1597341371
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1597341371
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1597341371
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1597341371
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1597341371
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1597341371
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1597341371
transform 1 0 15456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1597341371
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_160
timestamp 1597341371
transform 1 0 15824 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_160
timestamp 1597341371
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__SET_B
timestamp 1597341371
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__D
timestamp 1597341371
transform 1 0 15824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp 1597341371
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1597341371
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_167
timestamp 1597341371
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_163
timestamp 1597341371
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__CLK
timestamp 1597341371
transform 1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1597341371
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _201_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 16560 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _140_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 16652 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_4  _278_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 16376 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1597341371
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1597341371
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__D
timestamp 1597341371
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1597341371
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1597341371
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__B
timestamp 1597341371
transform 1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1597341371
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1597341371
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1597341371
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1597341371
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _146_
timestamp 1597341371
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1597341371
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1597341371
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1597341371
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_192
timestamp 1597341371
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1597341371
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1597341371
transform 1 0 18768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1597341371
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_198
timestamp 1597341371
transform 1 0 19320 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1597341371
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1597341371
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1597341371
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1597341371
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1597341371
transform 1 0 19136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1597341371
transform 1 0 19320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1597341371
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1597341371
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_203
timestamp 1597341371
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_208
timestamp 1597341371
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1597341371
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_200
timestamp 1597341371
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1597341371
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__D
timestamp 1597341371
transform 1 0 20056 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 1597341371
transform 1 0 19688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1597341371
transform 1 0 19596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1597341371
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1597341371
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1597341371
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1597341371
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_213
timestamp 1597341371
transform 1 0 20700 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_201
timestamp 1597341371
transform 1 0 19596 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1597341371
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1597341371
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1597341371
transform 1 0 22908 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1597341371
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1597341371
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1597341371
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1597341371
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1597341371
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1597341371
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1597341371
transform 1 0 21804 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1597341371
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1597341371
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1597341371
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1597341371
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1597341371
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1597341371
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1597341371
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1597341371
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1597341371
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1597341371
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_292
timestamp 1597341371
transform 1 0 27968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1597341371
transform 1 0 27600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_292
timestamp 1597341371
transform 1 0 27968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1597341371
transform -1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1597341371
transform -1 0 28336 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1597341371
transform -1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1597341371
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1597341371
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1597341371
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1597341371
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1597341371
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1597341371
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1597341371
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1597341371
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1597341371
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1597341371
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1597341371
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1597341371
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1597341371
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1597341371
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1597341371
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_62
timestamp 1597341371
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1597341371
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1597341371
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1597341371
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_74
timestamp 1597341371
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1597341371
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1597341371
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1597341371
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1597341371
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 1597341371
transform 1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A1
timestamp 1597341371
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1597341371
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_86
timestamp 1597341371
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1597341371
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 1597341371
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1597341371
transform 1 0 8740 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B1
timestamp 1597341371
transform 1 0 8096 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A2
timestamp 1597341371
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A1
timestamp 1597341371
transform 1 0 8832 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _205_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 8096 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp 1597341371
transform 1 0 10028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1597341371
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1597341371
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1597341371
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1597341371
transform 1 0 9200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__B1
timestamp 1597341371
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__RESET_B
timestamp 1597341371
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1597341371
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _291_
timestamp 1597341371
transform 1 0 9476 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1597341371
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1597341371
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1597341371
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1597341371
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1597341371
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1597341371
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1597341371
transform 1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A2
timestamp 1597341371
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1597341371
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _165_
timestamp 1597341371
transform 1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _204_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10488 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1597341371
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_130
timestamp 1597341371
transform 1 0 13064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1597341371
transform 1 0 12788 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1597341371
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__C
timestamp 1597341371
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _166_
timestamp 1597341371
transform 1 0 13340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_142
timestamp 1597341371
transform 1 0 14168 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1597341371
transform 1 0 13892 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1597341371
transform 1 0 13524 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_142
timestamp 1597341371
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1597341371
transform 1 0 13984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_147
timestamp 1597341371
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_146
timestamp 1597341371
transform 1 0 14536 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1597341371
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1597341371
transform 1 0 14444 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__B1
timestamp 1597341371
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1597341371
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_150
timestamp 1597341371
transform 1 0 14904 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__RESET_B
timestamp 1597341371
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1597341371
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1597341371
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1597341371
transform 1 0 15456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1597341371
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1597341371
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1597341371
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1597341371
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__CLK
timestamp 1597341371
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_162
timestamp 1597341371
transform 1 0 16008 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _173_
timestamp 1597341371
transform 1 0 16376 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _279_
timestamp 1597341371
transform 1 0 15824 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_4_183
timestamp 1597341371
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1597341371
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1597341371
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__B
timestamp 1597341371
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1597341371
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1597341371
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1597341371
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__C
timestamp 1597341371
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _200_
timestamp 1597341371
transform 1 0 18216 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp 1597341371
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_198
timestamp 1597341371
transform 1 0 19320 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1597341371
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1597341371
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A1
timestamp 1597341371
transform 1 0 19228 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1597341371
transform 1 0 19136 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_199
timestamp 1597341371
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1597341371
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1597341371
transform 1 0 19688 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1597341371
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1597341371
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1597341371
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1597341371
transform 1 0 20056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 1597341371
transform 1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1597341371
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1597341371
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_219
timestamp 1597341371
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1597341371
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1597341371
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__B
timestamp 1597341371
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A
timestamp 1597341371
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1597341371
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_223
timestamp 1597341371
transform 1 0 21620 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_212
timestamp 1597341371
transform 1 0 20608 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_247
timestamp 1597341371
transform 1 0 23828 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_235
timestamp 1597341371
transform 1 0 22724 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1597341371
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_236
timestamp 1597341371
transform 1 0 22816 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_224
timestamp 1597341371
transform 1 0 21712 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1597341371
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1597341371
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1597341371
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1597341371
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1597341371
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_292
timestamp 1597341371
transform 1 0 27968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1597341371
transform 1 0 27600 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1597341371
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1597341371
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1597341371
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1597341371
transform -1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1597341371
transform -1 0 28336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1597341371
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1597341371
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1597341371
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1597341371
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1597341371
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1597341371
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_44
timestamp 1597341371
transform 1 0 5152 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1597341371
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1597341371
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1597341371
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1597341371
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1597341371
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1597341371
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1597341371
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1597341371
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A3
timestamp 1597341371
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1597341371
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1597341371
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_62
timestamp 1597341371
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1597341371
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__D
timestamp 1597341371
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1597341371
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1597341371
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__RESET_B
timestamp 1597341371
transform 1 0 7084 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__CLK
timestamp 1597341371
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_67
timestamp 1597341371
transform 1 0 7268 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1597341371
transform 1 0 7268 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_71
timestamp 1597341371
transform 1 0 7636 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 1597341371
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_71
timestamp 1597341371
transform 1 0 7636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__B
timestamp 1597341371
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _272_
timestamp 1597341371
transform 1 0 7728 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1597341371
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_78
timestamp 1597341371
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B2
timestamp 1597341371
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B2
timestamp 1597341371
transform 1 0 8096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B1
timestamp 1597341371
transform 1 0 8556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1597341371
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_87
timestamp 1597341371
transform 1 0 9108 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_83
timestamp 1597341371
transform 1 0 8740 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1597341371
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_83
timestamp 1597341371
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B
timestamp 1597341371
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A2
timestamp 1597341371
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _148_
timestamp 1597341371
transform 1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1597341371
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_96
timestamp 1597341371
transform 1 0 9936 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1597341371
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A
timestamp 1597341371
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1597341371
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _274_
timestamp 1597341371
transform 1 0 9844 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_6_110
timestamp 1597341371
transform 1 0 11224 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_106
timestamp 1597341371
transform 1 0 10856 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1597341371
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__B1
timestamp 1597341371
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _196_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 11316 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1597341371
transform 1 0 12512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1597341371
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1597341371
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1597341371
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1597341371
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__D
timestamp 1597341371
transform 1 0 12328 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__D
timestamp 1597341371
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1597341371
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _169_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10304 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1597341371
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _178_
timestamp 1597341371
transform 1 0 12880 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _167_
timestamp 1597341371
transform 1 0 12604 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1597341371
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1597341371
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1597341371
transform 1 0 14260 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_138
timestamp 1597341371
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__B
timestamp 1597341371
transform 1 0 13616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B1
timestamp 1597341371
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A2
timestamp 1597341371
transform 1 0 13892 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1597341371
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1597341371
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1597341371
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1597341371
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__C1
timestamp 1597341371
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_160
timestamp 1597341371
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1597341371
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1597341371
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_160
timestamp 1597341371
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1597341371
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _179_
timestamp 1597341371
transform 1 0 14996 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _160_
timestamp 1597341371
transform 1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1597341371
transform 1 0 16192 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1597341371
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A1
timestamp 1597341371
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A2
timestamp 1597341371
transform 1 0 16008 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _269_
timestamp 1597341371
transform 1 0 16560 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _214_
timestamp 1597341371
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1597341371
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1597341371
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1597341371
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B1
timestamp 1597341371
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1597341371
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1597341371
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_187
timestamp 1597341371
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_184
timestamp 1597341371
transform 1 0 18032 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1597341371
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__D
timestamp 1597341371
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__CLK
timestamp 1597341371
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _222_
timestamp 1597341371
transform 1 0 18860 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _199_
timestamp 1597341371
transform 1 0 18216 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_195
timestamp 1597341371
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__B2
timestamp 1597341371
transform 1 0 19228 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_204
timestamp 1597341371
transform 1 0 19872 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_200
timestamp 1597341371
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_199
timestamp 1597341371
transform 1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__RESET_B
timestamp 1597341371
transform 1 0 19688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _216_
timestamp 1597341371
transform 1 0 19688 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1597341371
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1597341371
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1597341371
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B1
timestamp 1597341371
transform 1 0 20516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A2
timestamp 1597341371
transform 1 0 20240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1597341371
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_220
timestamp 1597341371
transform 1 0 21344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp 1597341371
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1597341371
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1597341371
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B
timestamp 1597341371
transform 1 0 21252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B2
timestamp 1597341371
transform 1 0 20884 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__RESET_B
timestamp 1597341371
transform 1 0 21528 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__D
timestamp 1597341371
transform 1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1597341371
transform 1 0 21620 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1597341371
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1597341371
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1597341371
transform 1 0 22264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__B1
timestamp 1597341371
transform 1 0 21896 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1597341371
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_237
timestamp 1597341371
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1597341371
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_244
timestamp 1597341371
transform 1 0 23552 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_232
timestamp 1597341371
transform 1 0 22448 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1597341371
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1597341371
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_268
timestamp 1597341371
transform 1 0 25760 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_256
timestamp 1597341371
transform 1 0 24656 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1597341371
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1597341371
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_292
timestamp 1597341371
transform 1 0 27968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1597341371
transform 1 0 27600 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1597341371
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1597341371
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1597341371
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1597341371
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1597341371
transform -1 0 28336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1597341371
transform -1 0 28336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1597341371
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1597341371
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1597341371
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1597341371
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1597341371
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1597341371
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1597341371
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1597341371
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1597341371
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 1597341371
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1597341371
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1597341371
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1597341371
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1597341371
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_56
timestamp 1597341371
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1597341371
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1597341371
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_53
timestamp 1597341371
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A2
timestamp 1597341371
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A1
timestamp 1597341371
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1597341371
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1597341371
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1597341371
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__B
timestamp 1597341371
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _293_
timestamp 1597341371
transform 1 0 7084 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__a32o_4  _276_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7268 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_8_84
timestamp 1597341371
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1597341371
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1597341371
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp 1597341371
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1597341371
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1597341371
transform 1 0 9200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A
timestamp 1597341371
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1597341371
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _171_
timestamp 1597341371
transform 1 0 10028 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _275_
timestamp 1597341371
transform 1 0 9936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_110
timestamp 1597341371
transform 1 0 11224 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp 1597341371
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1597341371
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1597341371
transform 1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__C
timestamp 1597341371
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1597341371
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__B
timestamp 1597341371
transform 1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__RESET_B
timestamp 1597341371
transform 1 0 11592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1597341371
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1597341371
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1597341371
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1597341371
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1597341371
transform 1 0 11960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__CLK
timestamp 1597341371
transform 1 0 11960 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1597341371
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1597341371
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _292_
timestamp 1597341371
transform 1 0 12328 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1597341371
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1597341371
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1597341371
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1597341371
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_137
timestamp 1597341371
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__B
timestamp 1597341371
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1597341371
transform 1 0 14260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1597341371
transform 1 0 14628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1597341371
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _197_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1597341371
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1597341371
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_156
timestamp 1597341371
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_150
timestamp 1597341371
transform 1 0 14904 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1597341371
transform 1 0 15456 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B
timestamp 1597341371
transform 1 0 15272 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1597341371
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_169
timestamp 1597341371
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1597341371
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1597341371
transform 1 0 16928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _180_
timestamp 1597341371
transform 1 0 16008 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _270_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15640 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp 1597341371
transform 1 0 17112 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_176
timestamp 1597341371
transform 1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__B
timestamp 1597341371
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A2
timestamp 1597341371
transform 1 0 17112 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1597341371
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1597341371
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A2
timestamp 1597341371
transform 1 0 17572 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1597341371
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _221_
timestamp 1597341371
transform 1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1597341371
transform 1 0 18032 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1597341371
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1597341371
transform 1 0 18216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1597341371
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_188
timestamp 1597341371
transform 1 0 18400 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__C
timestamp 1597341371
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _281_
timestamp 1597341371
transform 1 0 18768 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__o22a_4  _215_
timestamp 1597341371
transform 1 0 18768 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1597341371
transform 1 0 20056 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 1597341371
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 1597341371
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1597341371
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp 1597341371
transform 1 0 21344 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_215
timestamp 1597341371
transform 1 0 20884 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__CLK
timestamp 1597341371
transform 1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1597341371
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _218_
timestamp 1597341371
transform 1 0 21620 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _282_
timestamp 1597341371
transform 1 0 21160 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_8_245
timestamp 1597341371
transform 1 0 23644 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_241
timestamp 1597341371
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1597341371
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_236
timestamp 1597341371
transform 1 0 22816 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_232
timestamp 1597341371
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A1
timestamp 1597341371
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1597341371
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1597341371
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_269
timestamp 1597341371
transform 1 0 25852 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_257
timestamp 1597341371
transform 1 0 24748 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1597341371
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1597341371
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_292
timestamp 1597341371
transform 1 0 27968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1597341371
transform 1 0 27600 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1597341371
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1597341371
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1597341371
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1597341371
transform -1 0 28336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1597341371
transform -1 0 28336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1597341371
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1597341371
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1597341371
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1597341371
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1597341371
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1597341371
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1597341371
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1597341371
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1597341371
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1597341371
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1597341371
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1597341371
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_56
timestamp 1597341371
transform 1 0 6256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1597341371
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1597341371
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1597341371
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1597341371
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1597341371
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1597341371
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_68
timestamp 1597341371
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A2
timestamp 1597341371
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1597341371
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1597341371
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _273_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7544 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _271_
timestamp 1597341371
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1597341371
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1597341371
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1597341371
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__B1
timestamp 1597341371
transform 1 0 8556 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1597341371
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1597341371
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp 1597341371
transform 1 0 9108 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A1
timestamp 1597341371
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__B
timestamp 1597341371
transform 1 0 9016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1597341371
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _177_
timestamp 1597341371
transform 1 0 9384 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1597341371
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1597341371
transform 1 0 10212 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__B
timestamp 1597341371
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1597341371
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1597341371
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1597341371
transform 1 0 10580 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__C
timestamp 1597341371
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1597341371
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1597341371
transform 1 0 10672 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _185_
timestamp 1597341371
transform 1 0 10672 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_117
timestamp 1597341371
transform 1 0 11868 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1597341371
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1597341371
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1597341371
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 1597341371
transform 1 0 11592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1597341371
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1597341371
transform 1 0 11960 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1597341371
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1597341371
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1597341371
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__CLK
timestamp 1597341371
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__RESET_B
timestamp 1597341371
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1597341371
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1597341371
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1597341371
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1597341371
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1597341371
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__B1
timestamp 1597341371
transform 1 0 13432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__D
timestamp 1597341371
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _168_
timestamp 1597341371
transform 1 0 12604 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1597341371
transform 1 0 14720 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1597341371
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_145
timestamp 1597341371
transform 1 0 14444 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1597341371
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A1
timestamp 1597341371
transform 1 0 14260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1597341371
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B2
timestamp 1597341371
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1597341371
transform 1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _266_
timestamp 1597341371
transform 1 0 13248 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1597341371
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1597341371
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1597341371
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1597341371
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1597341371
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1597341371
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1597341371
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _209_
timestamp 1597341371
transform 1 0 15088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1597341371
transform 1 0 16652 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1597341371
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A2_N
timestamp 1597341371
transform 1 0 16468 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A1_N
timestamp 1597341371
transform 1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _184_
timestamp 1597341371
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _268_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15824 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_180
timestamp 1597341371
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_176
timestamp 1597341371
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1597341371
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1597341371
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1597341371
transform 1 0 17388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__RESET_B
timestamp 1597341371
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__D
timestamp 1597341371
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1597341371
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_188
timestamp 1597341371
transform 1 0 18400 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1597341371
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1597341371
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp 1597341371
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__B
timestamp 1597341371
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__D
timestamp 1597341371
transform 1 0 18308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _219_
timestamp 1597341371
transform 1 0 18676 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _207_
timestamp 1597341371
transform 1 0 18676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 1597341371
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_204
timestamp 1597341371
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1597341371
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_204
timestamp 1597341371
transform 1 0 19872 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1597341371
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1597341371
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1597341371
transform 1 0 19688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A3
timestamp 1597341371
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__B2
timestamp 1597341371
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1597341371
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1597341371
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1597341371
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1597341371
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _226_
timestamp 1597341371
transform 1 0 21068 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _223_
timestamp 1597341371
transform 1 0 20240 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1597341371
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_226
timestamp 1597341371
transform 1 0 21896 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B2
timestamp 1597341371
transform 1 0 22724 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B1
timestamp 1597341371
transform 1 0 21712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1597341371
transform 1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1597341371
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1597341371
transform 1 0 22908 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1597341371
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_243
timestamp 1597341371
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_231
timestamp 1597341371
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1597341371
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1597341371
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_255
timestamp 1597341371
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1597341371
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1597341371
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_292
timestamp 1597341371
transform 1 0 27968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_288
timestamp 1597341371
transform 1 0 27600 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1597341371
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1597341371
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1597341371
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1597341371
transform -1 0 28336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1597341371
transform -1 0 28336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1597341371
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1597341371
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1597341371
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1597341371
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1597341371
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1597341371
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1597341371
transform 1 0 5152 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1597341371
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1597341371
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1597341371
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1597341371
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1597341371
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1597341371
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1597341371
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1597341371
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 1597341371
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__B2
timestamp 1597341371
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1597341371
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1597341371
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1597341371
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1597341371
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A3
timestamp 1597341371
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1597341371
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1597341371
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _142_
timestamp 1597341371
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_74
timestamp 1597341371
transform 1 0 7912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_69
timestamp 1597341371
transform 1 0 7452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_72
timestamp 1597341371
transform 1 0 7728 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_68
timestamp 1597341371
transform 1 0 7360 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__B
timestamp 1597341371
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A1
timestamp 1597341371
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1597341371
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1597341371
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1597341371
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1597341371
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _192_
timestamp 1597341371
transform 1 0 8556 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _186_
timestamp 1597341371
transform 1 0 8188 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1597341371
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1597341371
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_94
timestamp 1597341371
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_88
timestamp 1597341371
transform 1 0 9200 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B
timestamp 1597341371
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__B1
timestamp 1597341371
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1597341371
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _208_
timestamp 1597341371
transform 1 0 9936 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _172_
timestamp 1597341371
transform 1 0 9844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1597341371
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1597341371
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_109
timestamp 1597341371
transform 1 0 11132 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1597341371
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1597341371
transform 1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__RESET_B
timestamp 1597341371
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_112
timestamp 1597341371
transform 1 0 11408 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1597341371
transform 1 0 11868 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B
timestamp 1597341371
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1597341371
transform 1 0 11960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _139_
timestamp 1597341371
transform 1 0 11960 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1597341371
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1597341371
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1597341371
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1597341371
transform 1 0 13524 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_131
timestamp 1597341371
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1597341371
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1597341371
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A2
timestamp 1597341371
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1597341371
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp 1597341371
transform 1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 1597341371
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1597341371
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1597341371
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1597341371
transform 1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1597341371
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1597341371
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _296_
timestamp 1597341371
transform 1 0 12972 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1597341371
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1597341371
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1597341371
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1597341371
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__B
timestamp 1597341371
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1597341371
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1597341371
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _213_
timestamp 1597341371
transform 1 0 15456 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1597341371
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1597341371
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_164
timestamp 1597341371
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1597341371
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1597341371
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__B1
timestamp 1597341371
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _182_
timestamp 1597341371
transform 1 0 16376 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_171
timestamp 1597341371
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1597341371
transform 1 0 16652 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1597341371
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1597341371
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1597341371
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__CLK
timestamp 1597341371
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1597341371
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _183_
timestamp 1597341371
transform 1 0 18216 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1597341371
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_198
timestamp 1597341371
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp 1597341371
transform 1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A2
timestamp 1597341371
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _280_
timestamp 1597341371
transform 1 0 17112 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1597341371
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_205
timestamp 1597341371
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1597341371
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1597341371
transform 1 0 20148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__B1
timestamp 1597341371
transform 1 0 19780 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1597341371
transform 1 0 19412 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1597341371
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1597341371
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1597341371
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_218
timestamp 1597341371
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A2
timestamp 1597341371
transform 1 0 21344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1597341371
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _227_
timestamp 1597341371
transform 1 0 21068 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__o32a_4  _212_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 19504 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_11_234
timestamp 1597341371
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_230
timestamp 1597341371
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_226
timestamp 1597341371
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A2_N
timestamp 1597341371
transform 1 0 22448 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1_N
timestamp 1597341371
transform 1 0 22080 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__B2
timestamp 1597341371
transform 1 0 21712 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_238
timestamp 1597341371
transform 1 0 23000 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__B1
timestamp 1597341371
transform 1 0 22816 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1597341371
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_245
timestamp 1597341371
transform 1 0 23644 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1597341371
transform 1 0 22540 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1597341371
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_269
timestamp 1597341371
transform 1 0 25852 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_257
timestamp 1597341371
transform 1 0 24748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1597341371
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1597341371
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_292
timestamp 1597341371
transform 1 0 27968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1597341371
transform 1 0 27600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1597341371
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1597341371
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1597341371
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1597341371
transform -1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1597341371
transform -1 0 28336 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1597341371
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1597341371
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1597341371
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1597341371
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1597341371
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1597341371
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1597341371
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1597341371
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1597341371
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1597341371
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1597341371
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1597341371
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1597341371
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1597341371
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1597341371
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1597341371
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1597341371
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1597341371
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__RESET_B
timestamp 1597341371
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1597341371
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1597341371
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1597341371
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__D
timestamp 1597341371
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__CLK
timestamp 1597341371
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _295_
timestamp 1597341371
transform 1 0 6716 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__a32o_4  _194_
timestamp 1597341371
transform 1 0 7728 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1597341371
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1597341371
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_89
timestamp 1597341371
transform 1 0 9292 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A1_N
timestamp 1597341371
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1597341371
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1597341371
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1597341371
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1597341371
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1597341371
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__B1
timestamp 1597341371
transform 1 0 10028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1597341371
transform 1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_99
timestamp 1597341371
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1597341371
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1597341371
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A2_N
timestamp 1597341371
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__CLK
timestamp 1597341371
transform 1 0 11316 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _170_
timestamp 1597341371
transform 1 0 10488 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1597341371
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1597341371
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1597341371
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1597341371
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__D
timestamp 1597341371
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1597341371
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _294_
timestamp 1597341371
transform 1 0 10856 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_14_129
timestamp 1597341371
transform 1 0 12972 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_128
timestamp 1597341371
transform 1 0 12880 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__RESET_B
timestamp 1597341371
transform 1 0 13340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1597341371
transform 1 0 12604 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1597341371
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1597341371
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1597341371
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1597341371
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__CLK
timestamp 1597341371
transform 1 0 14168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _261_
timestamp 1597341371
transform 1 0 13984 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp 1597341371
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1597341371
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1597341371
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1597341371
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__D
timestamp 1597341371
transform 1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1597341371
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1597341371
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A1
timestamp 1597341371
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1597341371
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1597341371
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A2
timestamp 1597341371
transform 1 0 15456 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B1
timestamp 1597341371
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_158
timestamp 1597341371
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_159
timestamp 1597341371
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__C1
timestamp 1597341371
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1_N
timestamp 1597341371
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_162
timestamp 1597341371
transform 1 0 16008 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1597341371
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1597341371
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1597341371
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A2_N
timestamp 1597341371
transform 1 0 16284 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1597341371
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _267_
timestamp 1597341371
transform 1 0 16376 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_182
timestamp 1597341371
transform 1 0 17848 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1597341371
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1597341371
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1597341371
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B1
timestamp 1597341371
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1597341371
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B2
timestamp 1597341371
transform 1 0 17112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1597341371
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1597341371
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp 1597341371
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1597341371
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1597341371
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_188
timestamp 1597341371
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1597341371
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A2
timestamp 1597341371
transform 1 0 18860 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__C
timestamp 1597341371
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _225_
timestamp 1597341371
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _220_
timestamp 1597341371
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1597341371
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1597341371
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__C1
timestamp 1597341371
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__B1
timestamp 1597341371
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1597341371
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_213
timestamp 1597341371
transform 1 0 20700 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1597341371
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__B
timestamp 1597341371
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1597341371
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__D
timestamp 1597341371
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1597341371
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp 1597341371
transform 1 0 20976 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1597341371
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_219
timestamp 1597341371
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A1
timestamp 1597341371
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1597341371
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_223
timestamp 1597341371
transform 1 0 21620 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_223
timestamp 1597341371
transform 1 0 21620 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1597341371
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_229
timestamp 1597341371
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__RESET_B
timestamp 1597341371
transform 1 0 22724 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__D
timestamp 1597341371
transform 1 0 22356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__CLK
timestamp 1597341371
transform 1 0 21988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_241
timestamp 1597341371
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_237
timestamp 1597341371
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__D
timestamp 1597341371
transform 1 0 23092 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1597341371
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1597341371
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _283_
timestamp 1597341371
transform 1 0 21988 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_14_262
timestamp 1597341371
transform 1 0 25208 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_250
timestamp 1597341371
transform 1 0 24104 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1597341371
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1597341371
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_292
timestamp 1597341371
transform 1 0 27968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1597341371
transform 1 0 27600 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1597341371
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1597341371
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1597341371
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1597341371
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1597341371
transform -1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1597341371
transform -1 0 28336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1597341371
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1597341371
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1597341371
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1597341371
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1597341371
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1597341371
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1597341371
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1597341371
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1597341371
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1597341371
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1597341371
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1597341371
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_68
timestamp 1597341371
transform 1 0 7360 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1597341371
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1597341371
transform 1 0 7820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1597341371
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1597341371
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1597341371
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1597341371
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _191_
timestamp 1597341371
transform 1 0 6992 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_83
timestamp 1597341371
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1597341371
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_76
timestamp 1597341371
transform 1 0 8096 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_79
timestamp 1597341371
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A1
timestamp 1597341371
transform 1 0 8188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A2
timestamp 1597341371
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B1
timestamp 1597341371
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__B2
timestamp 1597341371
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1597341371
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1597341371
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1597341371
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1597341371
transform 1 0 10028 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1597341371
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _189_
timestamp 1597341371
transform 1 0 8556 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_103
timestamp 1597341371
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_111
timestamp 1597341371
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1597341371
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1597341371
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A3
timestamp 1597341371
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A1
timestamp 1597341371
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B2
timestamp 1597341371
transform 1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B1
timestamp 1597341371
transform 1 0 10764 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1597341371
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1597341371
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1597341371
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_115
timestamp 1597341371
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A2
timestamp 1597341371
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1597341371
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1597341371
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1597341371
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _190_
timestamp 1597341371
transform 1 0 10764 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_16_126
timestamp 1597341371
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1597341371
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A2
timestamp 1597341371
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A1
timestamp 1597341371
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A1
timestamp 1597341371
transform 1 0 12880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1597341371
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1597341371
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B1
timestamp 1597341371
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1597341371
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1597341371
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B2
timestamp 1597341371
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A3
timestamp 1597341371
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_146
timestamp 1597341371
transform 1 0 14536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1597341371
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1597341371
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A2
timestamp 1597341371
transform 1 0 13984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__B1_N
timestamp 1597341371
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A1
timestamp 1597341371
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _288_
timestamp 1597341371
transform 1 0 13708 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1597341371
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1597341371
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1597341371
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1597341371
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1597341371
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_170
timestamp 1597341371
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1597341371
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1597341371
transform 1 0 16560 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__B1
timestamp 1597341371
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1597341371
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _224_
timestamp 1597341371
transform 1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _255_
timestamp 1597341371
transform 1 0 15456 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1597341371
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1597341371
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1597341371
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1597341371
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A1
timestamp 1597341371
transform 1 0 17388 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1597341371
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _210_
timestamp 1597341371
transform 1 0 18216 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_194
timestamp 1597341371
transform 1 0 18952 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_188
timestamp 1597341371
transform 1 0 18400 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1597341371
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1_N
timestamp 1597341371
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__B1
timestamp 1597341371
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _229_
timestamp 1597341371
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _252_
timestamp 1597341371
transform 1 0 17296 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1597341371
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1597341371
transform 1 0 19780 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1597341371
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__B
timestamp 1597341371
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A2_N
timestamp 1597341371
transform 1 0 19596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_219
timestamp 1597341371
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1597341371
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1597341371
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1597341371
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1597341371
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1597341371
transform 1 0 21620 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1597341371
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _259_
timestamp 1597341371
transform 1 0 21528 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _257_
timestamp 1597341371
transform 1 0 20148 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_16_235
timestamp 1597341371
transform 1 0 22724 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_231
timestamp 1597341371
transform 1 0 22356 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_233
timestamp 1597341371
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1597341371
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1597341371
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1597341371
transform 1 0 22724 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A2
timestamp 1597341371
transform 1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__B2
timestamp 1597341371
transform 1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__C
timestamp 1597341371
transform 1 0 22540 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1597341371
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_237
timestamp 1597341371
transform 1 0 22908 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A1
timestamp 1597341371
transform 1 0 22908 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1597341371
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1597341371
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1597341371
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1597341371
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1597341371
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1597341371
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1597341371
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_292
timestamp 1597341371
transform 1 0 27968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_288
timestamp 1597341371
transform 1 0 27600 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1597341371
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1597341371
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1597341371
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1597341371
transform -1 0 28336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1597341371
transform -1 0 28336 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1597341371
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1597341371
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1597341371
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1597341371
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1597341371
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1597341371
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1597341371
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1597341371
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1597341371
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1597341371
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1597341371
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1597341371
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_68
timestamp 1597341371
transform 1 0 7360 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1597341371
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_74
timestamp 1597341371
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1597341371
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1597341371
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1597341371
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1597341371
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1597341371
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_76
timestamp 1597341371
transform 1 0 8096 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_83
timestamp 1597341371
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_79
timestamp 1597341371
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1597341371
transform 1 0 9016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__B
timestamp 1597341371
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1597341371
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _187_
timestamp 1597341371
transform 1 0 8188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1597341371
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_97
timestamp 1597341371
transform 1 0 10028 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1597341371
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1597341371
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _193_
timestamp 1597341371
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1597341371
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1597341371
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1597341371
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1597341371
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__B1
timestamp 1597341371
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1597341371
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__RESET_B
timestamp 1597341371
transform 1 0 10580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__D
timestamp 1597341371
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp 1597341371
transform 1 0 11316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1597341371
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1597341371
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1597341371
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__CLK
timestamp 1597341371
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1597341371
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _287_
timestamp 1597341371
transform 1 0 11500 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1597341371
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_132
timestamp 1597341371
transform 1 0 13248 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_128
timestamp 1597341371
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1597341371
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A1
timestamp 1597341371
transform 1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _164_
timestamp 1597341371
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_148
timestamp 1597341371
transform 1 0 14720 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1597341371
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1597341371
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1597341371
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1597341371
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__C
timestamp 1597341371
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__D
timestamp 1597341371
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A3
timestamp 1597341371
transform 1 0 14168 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__B1
timestamp 1597341371
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _256_
timestamp 1597341371
transform 1 0 14352 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1597341371
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1597341371
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1597341371
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1597341371
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1597341371
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1597341371
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 1597341371
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A2
timestamp 1597341371
transform 1 0 16468 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1597341371
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B1
timestamp 1597341371
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _211_
timestamp 1597341371
transform 1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_4  _254_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15456 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1597341371
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1597341371
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1597341371
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__B
timestamp 1597341371
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1597341371
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1597341371
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1597341371
transform 1 0 18216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B
timestamp 1597341371
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1597341371
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _240_
timestamp 1597341371
transform 1 0 17388 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_18_188
timestamp 1597341371
transform 1 0 18400 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1597341371
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _246_
timestamp 1597341371
transform 1 0 18768 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _258_
timestamp 1597341371
transform 1 0 18768 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1597341371
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1597341371
transform 1 0 19780 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_199
timestamp 1597341371
transform 1 0 19412 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1597341371
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__B1
timestamp 1597341371
transform 1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 1597341371
transform 1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1597341371
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1597341371
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_212
timestamp 1597341371
transform 1 0 20608 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B
timestamp 1597341371
transform 1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1597341371
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _263_
timestamp 1597341371
transform 1 0 20976 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _198_
timestamp 1597341371
transform 1 0 21068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_220
timestamp 1597341371
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1597341371
transform 1 0 21528 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_224
timestamp 1597341371
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1597341371
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_229
timestamp 1597341371
transform 1 0 22172 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1597341371
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__B1
timestamp 1597341371
transform 1 0 22724 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A2
timestamp 1597341371
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A2
timestamp 1597341371
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_246
timestamp 1597341371
transform 1 0 23736 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_242
timestamp 1597341371
transform 1 0 23368 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1597341371
transform 1 0 23000 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_241
timestamp 1597341371
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_237
timestamp 1597341371
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1597341371
transform 1 0 23092 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__B
timestamp 1597341371
transform 1 0 23184 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1597341371
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1597341371
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _265_
timestamp 1597341371
transform 1 0 21896 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1597341371
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_269
timestamp 1597341371
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1597341371
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_292
timestamp 1597341371
transform 1 0 27968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1597341371
transform 1 0 27600 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1597341371
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1597341371
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1597341371
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1597341371
transform -1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1597341371
transform -1 0 28336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1597341371
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1597341371
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1597341371
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1597341371
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1597341371
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1597341371
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1597341371
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1597341371
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1597341371
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1597341371
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1597341371
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1597341371
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1597341371
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1597341371
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_74
timestamp 1597341371
transform 1 0 7912 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1597341371
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1597341371
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1597341371
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1597341371
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1597341371
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1597341371
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1597341371
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_80
timestamp 1597341371
transform 1 0 8464 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_91
timestamp 1597341371
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1597341371
transform 1 0 8740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1597341371
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _176_
timestamp 1597341371
transform 1 0 8648 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_105
timestamp 1597341371
transform 1 0 10764 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1597341371
transform 1 0 10580 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1597341371
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_111
timestamp 1597341371
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1597341371
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_111
timestamp 1597341371
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__C
timestamp 1597341371
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__B
timestamp 1597341371
transform 1 0 11592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1597341371
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1597341371
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1597341371
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1597341371
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1597341371
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__B2
timestamp 1597341371
transform 1 0 11960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B2
timestamp 1597341371
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A1
timestamp 1597341371
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1597341371
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1597341371
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_126
timestamp 1597341371
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__B1
timestamp 1597341371
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1597341371
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1597341371
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_146
timestamp 1597341371
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1597341371
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A2
timestamp 1597341371
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A2
timestamp 1597341371
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A1
timestamp 1597341371
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _251_
timestamp 1597341371
transform 1 0 12604 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_4  _250_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 13248 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1597341371
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_161
timestamp 1597341371
transform 1 0 15916 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1597341371
transform 1 0 15548 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_154
timestamp 1597341371
transform 1 0 15272 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1597341371
transform 1 0 14904 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__B
timestamp 1597341371
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1597341371
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _262_
timestamp 1597341371
transform 1 0 15456 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_171
timestamp 1597341371
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_165
timestamp 1597341371
transform 1 0 16284 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__B
timestamp 1597341371
transform 1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _238_
timestamp 1597341371
transform 1 0 17020 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _248_
timestamp 1597341371
transform 1 0 16008 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1597341371
transform 1 0 17664 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1597341371
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1597341371
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1597341371
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1597341371
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_187
timestamp 1597341371
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_184
timestamp 1597341371
transform 1 0 18032 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1597341371
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1597341371
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B2
timestamp 1597341371
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _237_
timestamp 1597341371
transform 1 0 18216 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _233_
timestamp 1597341371
transform 1 0 18492 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1597341371
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1597341371
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1597341371
transform 1 0 19044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp 1597341371
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_202
timestamp 1597341371
transform 1 0 19688 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 1597341371
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1597341371
transform 1 0 19412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1597341371
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 1597341371
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B1
timestamp 1597341371
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_220
timestamp 1597341371
transform 1 0 21344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1597341371
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1597341371
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1597341371
transform 1 0 21344 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_216
timestamp 1597341371
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__C
timestamp 1597341371
transform 1 0 21528 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1597341371
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1597341371
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _217_
timestamp 1597341371
transform 1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _260_
timestamp 1597341371
transform 1 0 19872 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_233
timestamp 1597341371
transform 1 0 22540 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _264_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 21712 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_244
timestamp 1597341371
transform 1 0 23552 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_236
timestamp 1597341371
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1597341371
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1597341371
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 1597341371
transform 1 0 23092 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_AMUX2_3V_I1
timestamp 1597341371
transform 1 0 23644 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_AMUX2_3V_select
timestamp 1597341371
transform 1 0 23184 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1597341371
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_247
timestamp 1597341371
transform 1 0 23828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_224
timestamp 1597341371
transform 1 0 21712 0 -1 13600
box -38 -48 1142 592
use AMUX2_3V  AMUX2_3V
timestamp 1598265745
transform 1 0 23828 0 1 11968
box 0 0 1812 1088
use sky130_fd_sc_hd__decap_4  FILLER_20_271
timestamp 1597341371
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_259
timestamp 1597341371
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_267
timestamp 1597341371
transform 1 0 25668 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_292
timestamp 1597341371
transform 1 0 27968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_288
timestamp 1597341371
transform 1 0 27600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1597341371
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_291
timestamp 1597341371
transform 1 0 27876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_279
timestamp 1597341371
transform 1 0 26772 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1597341371
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1597341371
transform -1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1597341371
transform -1 0 28336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1597341371
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1597341371
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1597341371
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1597341371
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1597341371
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1597341371
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1597341371
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1597341371
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1597341371
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1597341371
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1597341371
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1597341371
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1597341371
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1597341371
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_74
timestamp 1597341371
transform 1 0 7912 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1597341371
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1597341371
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1597341371
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1597341371
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1597341371
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1597341371
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1597341371
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1597341371
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1597341371
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1597341371
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _175_
timestamp 1597341371
transform 1 0 8740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_105
timestamp 1597341371
transform 1 0 10764 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_113
timestamp 1597341371
transform 1 0 11500 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1597341371
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1597341371
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1597341371
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B1
timestamp 1597341371
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A2
timestamp 1597341371
transform 1 0 11592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_122
timestamp 1597341371
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_118
timestamp 1597341371
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1597341371
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1597341371
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A3
timestamp 1597341371
transform 1 0 11960 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__D
timestamp 1597341371
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__CLK
timestamp 1597341371
transform 1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1597341371
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_126
timestamp 1597341371
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 1597341371
transform 1 0 13156 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1597341371
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 1597341371
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__RESET_B
timestamp 1597341371
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1597341371
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1597341371
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1597341371
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1597341371
transform 1 0 14628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _247_
timestamp 1597341371
transform 1 0 12880 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_4  _245_
timestamp 1597341371
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1597341371
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_153
timestamp 1597341371
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__C
timestamp 1597341371
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1597341371
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _253_
timestamp 1597341371
transform 1 0 15456 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _249_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15364 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_165
timestamp 1597341371
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_168
timestamp 1597341371
transform 1 0 16560 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_164
timestamp 1597341371
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__B
timestamp 1597341371
transform 1 0 16468 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1597341371
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_169
timestamp 1597341371
transform 1 0 16652 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1597341371
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _239_
timestamp 1597341371
transform 1 0 16928 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_186
timestamp 1597341371
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_181
timestamp 1597341371
transform 1 0 17756 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_184
timestamp 1597341371
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1597341371
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_178
timestamp 1597341371
transform 1 0 17480 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1597341371
transform 1 0 17112 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A2_N
timestamp 1597341371
transform 1 0 18032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A2
timestamp 1597341371
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1597341371
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1597341371
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_189
timestamp 1597341371
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1597341371
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A1
timestamp 1597341371
transform 1 0 18308 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _234_
timestamp 1597341371
transform 1 0 18676 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _230_
timestamp 1597341371
transform 1 0 18768 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1597341371
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_205
timestamp 1597341371
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1_N
timestamp 1597341371
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B2
timestamp 1597341371
transform 1 0 20148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1597341371
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1597341371
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_213
timestamp 1597341371
transform 1 0 20700 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1597341371
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A2
timestamp 1597341371
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__D
timestamp 1597341371
transform 1 0 21068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1597341371
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _231_
timestamp 1597341371
transform 1 0 20976 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_223
timestamp 1597341371
transform 1 0 21620 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1597341371
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1597341371
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_233
timestamp 1597341371
transform 1 0 22540 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_225
timestamp 1597341371
transform 1 0 21804 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__D
timestamp 1597341371
transform 1 0 22724 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__CLK
timestamp 1597341371
transform 1 0 22356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_241
timestamp 1597341371
transform 1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_237
timestamp 1597341371
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__RESET_B
timestamp 1597341371
transform 1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1597341371
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1597341371
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _297_
timestamp 1597341371
transform 1 0 22356 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1597341371
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_254
timestamp 1597341371
transform 1 0 24472 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1597341371
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1597341371
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_292
timestamp 1597341371
transform 1 0 27968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1597341371
transform 1 0 27600 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1597341371
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1597341371
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1597341371
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1597341371
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1597341371
transform -1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1597341371
transform -1 0 28336 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1597341371
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1597341371
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1597341371
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1597341371
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1597341371
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1597341371
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1597341371
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1597341371
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1597341371
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1597341371
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1597341371
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1597341371
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1597341371
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1597341371
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1597341371
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1597341371
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1597341371
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1597341371
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1597341371
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1597341371
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1597341371
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1597341371
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1597341371
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1597341371
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_117
timestamp 1597341371
transform 1 0 11868 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1597341371
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1597341371
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1597341371
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_110
timestamp 1597341371
transform 1 0 11224 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1597341371
transform 1 0 11960 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1597341371
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_136
timestamp 1597341371
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_130
timestamp 1597341371
transform 1 0 13064 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1597341371
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__B
timestamp 1597341371
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _154_
timestamp 1597341371
transform 1 0 12788 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1597341371
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1597341371
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1597341371
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__CLK
timestamp 1597341371
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _242_
timestamp 1597341371
transform 1 0 13800 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  _286_
timestamp 1597341371
transform 1 0 12604 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1597341371
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_152
timestamp 1597341371
transform 1 0 15088 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__D
timestamp 1597341371
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1597341371
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _244_
timestamp 1597341371
transform 1 0 15364 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _236_
timestamp 1597341371
transform 1 0 15456 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_165
timestamp 1597341371
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_168
timestamp 1597341371
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_164
timestamp 1597341371
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1597341371
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B2
timestamp 1597341371
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_173
timestamp 1597341371
transform 1 0 17020 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_169
timestamp 1597341371
transform 1 0 16652 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1597341371
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B1
timestamp 1597341371
transform 1 0 16744 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1597341371
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1597341371
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_176
timestamp 1597341371
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A2
timestamp 1597341371
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1597341371
transform 1 0 17112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1597341371
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1597341371
transform 1 0 18400 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_194
timestamp 1597341371
transform 1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_190
timestamp 1597341371
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1597341371
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B1
timestamp 1597341371
transform 1 0 18768 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _232_
timestamp 1597341371
transform 1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _241_
timestamp 1597341371
transform 1 0 17112 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__a2bb2o_4  _235_
timestamp 1597341371
transform 1 0 19228 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_207
timestamp 1597341371
transform 1 0 20148 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1597341371
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1597341371
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1597341371
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B2
timestamp 1597341371
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1597341371
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1597341371
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_217
timestamp 1597341371
transform 1 0 21068 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1597341371
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__CLK
timestamp 1597341371
transform 1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1597341371
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1597341371
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _284_
timestamp 1597341371
transform 1 0 21068 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_24_240
timestamp 1597341371
transform 1 0 23184 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1597341371
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1597341371
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_228
timestamp 1597341371
transform 1 0 22080 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1597341371
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__RESET_B
timestamp 1597341371
transform 1 0 21896 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1597341371
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1597341371
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_264
timestamp 1597341371
transform 1 0 25392 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_252
timestamp 1597341371
transform 1 0 24288 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1597341371
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1597341371
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1597341371
transform 1 0 27968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_288
timestamp 1597341371
transform 1 0 27600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1597341371
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1597341371
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1597341371
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1597341371
transform -1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1597341371
transform -1 0 28336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1597341371
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1597341371
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1597341371
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1597341371
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1597341371
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1597341371
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1597341371
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1597341371
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1597341371
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1597341371
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1597341371
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1597341371
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1597341371
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1597341371
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1597341371
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1597341371
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1597341371
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1597341371
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1597341371
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1597341371
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1597341371
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1597341371
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1597341371
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1597341371
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1597341371
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1597341371
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1597341371
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1597341371
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1597341371
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1597341371
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1597341371
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1597341371
transform 1 0 14076 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1597341371
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1597341371
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1597341371
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__RESET_B
timestamp 1597341371
transform 1 0 14076 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1597341371
transform 1 0 14168 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1597341371
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _285_
timestamp 1597341371
transform 1 0 14444 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_26_158
timestamp 1597341371
transform 1 0 15640 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1597341371
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1597341371
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1597341371
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1597341371
transform 1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1597341371
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1597341371
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _243_
timestamp 1597341371
transform 1 0 15916 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1597341371
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 1597341371
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B1
timestamp 1597341371
transform 1 0 17112 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1597341371
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1597341371
transform 1 0 19136 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _228_
timestamp 1597341371
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_198
timestamp 1597341371
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_186
timestamp 1597341371
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_174
timestamp 1597341371
transform 1 0 17112 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1597341371
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1597341371
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1597341371
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_218
timestamp 1597341371
transform 1 0 21160 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_206
timestamp 1597341371
transform 1 0 20056 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1597341371
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1597341371
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1597341371
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1597341371
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_242
timestamp 1597341371
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_230
timestamp 1597341371
transform 1 0 22264 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1597341371
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1597341371
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1597341371
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1597341371
transform 1 0 25852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1597341371
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_292
timestamp 1597341371
transform 1 0 27968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1597341371
transform 1 0 27600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1597341371
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1597341371
transform 1 0 26956 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1597341371
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1597341371
transform -1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1597341371
transform -1 0 28336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1597341371
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1597341371
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1597341371
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1597341371
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1597341371
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1597341371
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1597341371
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1597341371
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1597341371
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1597341371
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1597341371
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1597341371
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1597341371
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1597341371
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1597341371
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1597341371
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1597341371
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1597341371
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1597341371
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1597341371
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1597341371
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1597341371
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1597341371
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1597341371
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1597341371
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1597341371
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1597341371
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1597341371
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1597341371
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1597341371
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1597341371
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1597341371
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1597341371
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1597341371
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1597341371
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1597341371
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1597341371
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1597341371
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1597341371
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1597341371
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1597341371
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1597341371
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1597341371
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1597341371
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1597341371
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1597341371
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1597341371
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1597341371
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1597341371
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1597341371
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1597341371
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1597341371
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1597341371
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1597341371
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1597341371
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1597341371
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1597341371
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_292
timestamp 1597341371
transform 1 0 27968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1597341371
transform 1 0 27600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1597341371
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1597341371
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1597341371
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1597341371
transform -1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1597341371
transform -1 0 28336 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1597341371
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1597341371
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1597341371
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1597341371
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1597341371
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1597341371
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1597341371
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1597341371
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1597341371
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1597341371
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1597341371
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1597341371
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1597341371
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1597341371
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1597341371
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1597341371
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1597341371
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1597341371
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1597341371
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1597341371
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1597341371
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1597341371
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1597341371
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1597341371
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1597341371
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1597341371
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1597341371
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1597341371
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1597341371
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1597341371
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1597341371
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1597341371
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1597341371
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1597341371
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1597341371
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1597341371
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1597341371
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1597341371
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1597341371
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1597341371
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1597341371
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1597341371
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1597341371
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1597341371
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1597341371
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1597341371
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1597341371
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1597341371
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1597341371
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1597341371
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1597341371
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1597341371
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1597341371
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1597341371
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1597341371
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1597341371
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1597341371
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_292
timestamp 1597341371
transform 1 0 27968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_288
timestamp 1597341371
transform 1 0 27600 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1597341371
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1597341371
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1597341371
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1597341371
transform -1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1597341371
transform -1 0 28336 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1597341371
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1597341371
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1597341371
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1597341371
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1597341371
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1597341371
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1597341371
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1597341371
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1597341371
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1597341371
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1597341371
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1597341371
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1597341371
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1597341371
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1597341371
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1597341371
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1597341371
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1597341371
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1597341371
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1597341371
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1597341371
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1597341371
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1597341371
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1597341371
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1597341371
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1597341371
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1597341371
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1597341371
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1597341371
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1597341371
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1597341371
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1597341371
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1597341371
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1597341371
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1597341371
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1597341371
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1597341371
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1597341371
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1597341371
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1597341371
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1597341371
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1597341371
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1597341371
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1597341371
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1597341371
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1597341371
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1597341371
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1597341371
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1597341371
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1597341371
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1597341371
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1597341371
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1597341371
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1597341371
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1597341371
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1597341371
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1597341371
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_292
timestamp 1597341371
transform 1 0 27968 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1597341371
transform 1 0 27600 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1597341371
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1597341371
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1597341371
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1597341371
transform -1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1597341371
transform -1 0 28336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1597341371
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1597341371
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1597341371
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1597341371
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1597341371
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1597341371
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1597341371
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1597341371
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1597341371
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1597341371
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1597341371
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1597341371
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1597341371
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1597341371
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1597341371
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1597341371
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1597341371
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1597341371
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1597341371
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1597341371
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1597341371
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1597341371
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1597341371
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1597341371
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1597341371
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1597341371
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1597341371
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1597341371
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1597341371
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1597341371
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1597341371
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1597341371
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1597341371
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1597341371
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1597341371
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1597341371
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1597341371
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1597341371
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1597341371
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1597341371
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1597341371
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1597341371
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1597341371
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1597341371
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1597341371
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1597341371
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1597341371
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1597341371
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1597341371
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1597341371
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1597341371
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1597341371
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1597341371
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1597341371
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1597341371
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1597341371
transform 1 0 25852 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1597341371
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_292
timestamp 1597341371
transform 1 0 27968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1597341371
transform 1 0 27600 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1597341371
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1597341371
transform 1 0 26956 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1597341371
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1597341371
transform -1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1597341371
transform -1 0 28336 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1597341371
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1597341371
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1597341371
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1597341371
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1597341371
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1597341371
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1597341371
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1597341371
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1597341371
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1597341371
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1597341371
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1597341371
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1597341371
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1597341371
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1597341371
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1597341371
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1597341371
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1597341371
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1597341371
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1597341371
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1597341371
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1597341371
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1597341371
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1597341371
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1597341371
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1597341371
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1597341371
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1597341371
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1597341371
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1597341371
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1597341371
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1597341371
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1597341371
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1597341371
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1597341371
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1597341371
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1597341371
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1597341371
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1597341371
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1597341371
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1597341371
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1597341371
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1597341371
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1597341371
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1597341371
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1597341371
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1597341371
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1597341371
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1597341371
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1597341371
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1597341371
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1597341371
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1597341371
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1597341371
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1597341371
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_269
timestamp 1597341371
transform 1 0 25852 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1597341371
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_292
timestamp 1597341371
transform 1 0 27968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1597341371
transform 1 0 27600 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1597341371
transform 1 0 26496 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1597341371
transform 1 0 26956 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1597341371
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1597341371
transform -1 0 28336 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1597341371
transform -1 0 28336 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1597341371
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1597341371
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1597341371
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1597341371
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1597341371
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1597341371
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1597341371
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1597341371
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1597341371
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1597341371
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1597341371
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1597341371
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1597341371
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1597341371
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1597341371
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1597341371
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1597341371
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1597341371
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1597341371
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1597341371
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1597341371
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1597341371
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1597341371
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1597341371
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1597341371
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1597341371
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1597341371
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1597341371
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1597341371
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1597341371
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1597341371
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1597341371
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1597341371
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1597341371
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1597341371
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1597341371
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1597341371
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1597341371
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1597341371
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1597341371
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1597341371
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1597341371
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1597341371
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1597341371
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1597341371
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1597341371
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1597341371
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1597341371
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1597341371
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1597341371
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1597341371
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1597341371
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1597341371
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1597341371
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1597341371
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_269
timestamp 1597341371
transform 1 0 25852 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1597341371
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_292
timestamp 1597341371
transform 1 0 27968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1597341371
transform 1 0 27600 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1597341371
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1597341371
transform 1 0 26956 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1597341371
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1597341371
transform -1 0 28336 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1597341371
transform -1 0 28336 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1597341371
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1597341371
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1597341371
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1597341371
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1597341371
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1597341371
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1597341371
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1597341371
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1597341371
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1597341371
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1597341371
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1597341371
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1597341371
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1597341371
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1597341371
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1597341371
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1597341371
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1597341371
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1597341371
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1597341371
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1597341371
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1597341371
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1597341371
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1597341371
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1597341371
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1597341371
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1597341371
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1597341371
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1597341371
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1597341371
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1597341371
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1597341371
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1597341371
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1597341371
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1597341371
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1597341371
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1597341371
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1597341371
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1597341371
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1597341371
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1597341371
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1597341371
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1597341371
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1597341371
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1597341371
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1597341371
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1597341371
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1597341371
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1597341371
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1597341371
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1597341371
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1597341371
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1597341371
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1597341371
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1597341371
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1597341371
transform 1 0 25852 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1597341371
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_292
timestamp 1597341371
transform 1 0 27968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1597341371
transform 1 0 27600 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1597341371
transform 1 0 26496 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1597341371
transform 1 0 26956 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1597341371
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1597341371
transform -1 0 28336 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1597341371
transform -1 0 28336 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1597341371
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1597341371
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1597341371
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1597341371
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1597341371
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1597341371
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1597341371
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1597341371
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1597341371
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1597341371
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1597341371
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1597341371
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1597341371
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1597341371
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1597341371
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1597341371
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1597341371
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1597341371
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1597341371
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1597341371
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_80
timestamp 1597341371
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1597341371
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1597341371
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1597341371
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_117
timestamp 1597341371
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1597341371
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1597341371
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1597341371
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1597341371
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1597341371
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1597341371
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1597341371
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1597341371
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_166
timestamp 1597341371
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1597341371
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1597341371
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1597341371
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1597341371
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_190
timestamp 1597341371
transform 1 0 18584 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_178
timestamp 1597341371
transform 1 0 17480 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1597341371
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1597341371
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1597341371
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1597341371
transform 1 0 20884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_202
timestamp 1597341371
transform 1 0 19688 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1597341371
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1597341371
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1597341371
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1597341371
transform 1 0 23092 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1597341371
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1597341371
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1597341371
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1597341371
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1597341371
transform 1 0 25300 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_251
timestamp 1597341371
transform 1 0 24196 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_269
timestamp 1597341371
transform 1 0 25852 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1597341371
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_292
timestamp 1597341371
transform 1 0 27968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_288
timestamp 1597341371
transform 1 0 27600 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1597341371
transform 1 0 26496 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1597341371
transform 1 0 26956 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1597341371
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1597341371
transform -1 0 28336 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1597341371
transform -1 0 28336 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1597341371
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1597341371
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1597341371
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1597341371
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1597341371
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1597341371
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1597341371
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1597341371
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1597341371
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1597341371
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1597341371
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1597341371
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1597341371
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_56
timestamp 1597341371
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_74
timestamp 1597341371
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1597341371
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1597341371
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_51
timestamp 1597341371
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1597341371
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1597341371
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_80
timestamp 1597341371
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_98
timestamp 1597341371
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_86
timestamp 1597341371
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1597341371
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1597341371
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1597341371
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1597341371
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_110
timestamp 1597341371
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1597341371
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1597341371
transform 1 0 14076 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1597341371
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_147
timestamp 1597341371
transform 1 0 14628 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1597341371
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_166
timestamp 1597341371
transform 1 0 16376 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1597341371
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_171
timestamp 1597341371
transform 1 0 16836 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_159
timestamp 1597341371
transform 1 0 15732 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1597341371
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_190
timestamp 1597341371
transform 1 0 18584 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_178
timestamp 1597341371
transform 1 0 17480 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1597341371
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1597341371
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1597341371
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1597341371
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_202
timestamp 1597341371
transform 1 0 19688 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1597341371
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1597341371
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1597341371
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_239
timestamp 1597341371
transform 1 0 23092 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1597341371
transform 1 0 21988 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1597341371
transform 1 0 23644 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1597341371
transform 1 0 22448 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1597341371
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_263
timestamp 1597341371
transform 1 0 25300 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_251
timestamp 1597341371
transform 1 0 24196 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_269
timestamp 1597341371
transform 1 0 25852 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1597341371
transform 1 0 24748 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_292
timestamp 1597341371
transform 1 0 27968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1597341371
transform 1 0 27600 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_276
timestamp 1597341371
transform 1 0 26496 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1597341371
transform 1 0 26956 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1597341371
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1597341371
transform -1 0 28336 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1597341371
transform -1 0 28336 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1597341371
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1597341371
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1597341371
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1597341371
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1597341371
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1597341371
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1597341371
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1597341371
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1597341371
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1597341371
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1597341371
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1597341371
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1597341371
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1597341371
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_74
timestamp 1597341371
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_62
timestamp 1597341371
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1597341371
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_51
timestamp 1597341371
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1597341371
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1597341371
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_80
timestamp 1597341371
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_98
timestamp 1597341371
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_86
timestamp 1597341371
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1597341371
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1597341371
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1597341371
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1597341371
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_110
timestamp 1597341371
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1597341371
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1597341371
transform 1 0 14076 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1597341371
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_147
timestamp 1597341371
transform 1 0 14628 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_135
timestamp 1597341371
transform 1 0 13524 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_166
timestamp 1597341371
transform 1 0 16376 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_154
timestamp 1597341371
transform 1 0 15272 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1597341371
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_159
timestamp 1597341371
transform 1 0 15732 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1597341371
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_190
timestamp 1597341371
transform 1 0 18584 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_178
timestamp 1597341371
transform 1 0 17480 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1597341371
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1597341371
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1597341371
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1597341371
transform 1 0 20884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_202
timestamp 1597341371
transform 1 0 19688 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_220
timestamp 1597341371
transform 1 0 21344 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1597341371
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1597341371
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_248
timestamp 1597341371
transform 1 0 23920 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_227
timestamp 1597341371
transform 1 0 21988 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1597341371
transform 1 0 23644 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_241
timestamp 1597341371
transform 1 0 23276 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_238
timestamp 1597341371
transform 1 0 23000 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_232
timestamp 1597341371
transform 1 0 22448 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1597341371
transform 1 0 23092 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1597341371
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _277_
timestamp 1597341371
transform 1 0 23092 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_46_272
timestamp 1597341371
transform 1 0 26128 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_260
timestamp 1597341371
transform 1 0 25024 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_269
timestamp 1597341371
transform 1 0 25852 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_257
timestamp 1597341371
transform 1 0 24748 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_292
timestamp 1597341371
transform 1 0 27968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_288
timestamp 1597341371
transform 1 0 27600 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_276
timestamp 1597341371
transform 1 0 26496 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1597341371
transform 1 0 26956 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1597341371
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1597341371
transform -1 0 28336 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1597341371
transform -1 0 28336 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1597341371
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1597341371
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1597341371
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1597341371
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1597341371
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1597341371
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1597341371
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1597341371
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1597341371
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1597341371
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1597341371
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1597341371
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1597341371
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1597341371
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_74
timestamp 1597341371
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1597341371
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1597341371
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1597341371
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1597341371
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1597341371
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1597341371
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_98
timestamp 1597341371
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_86
timestamp 1597341371
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1597341371
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1597341371
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1597341371
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1597341371
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_110
timestamp 1597341371
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1597341371
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1597341371
transform 1 0 14076 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1597341371
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1597341371
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_135
timestamp 1597341371
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1597341371
transform 1 0 16376 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1597341371
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_171
timestamp 1597341371
transform 1 0 16836 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1597341371
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1597341371
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_190
timestamp 1597341371
transform 1 0 18584 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1597341371
transform 1 0 17480 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1597341371
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1597341371
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1597341371
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1597341371
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_202
timestamp 1597341371
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_220
timestamp 1597341371
transform 1 0 21344 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1597341371
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1597341371
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1597341371
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1597341371
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_245
timestamp 1597341371
transform 1 0 23644 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_232
timestamp 1597341371
transform 1 0 22448 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1597341371
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_263
timestamp 1597341371
transform 1 0 25300 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_251
timestamp 1597341371
transform 1 0 24196 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_269
timestamp 1597341371
transform 1 0 25852 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_257
timestamp 1597341371
transform 1 0 24748 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_292
timestamp 1597341371
transform 1 0 27968 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_288
timestamp 1597341371
transform 1 0 27600 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_276
timestamp 1597341371
transform 1 0 26496 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1597341371
transform 1 0 26956 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1597341371
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1597341371
transform -1 0 28336 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1597341371
transform -1 0 28336 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1597341371
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1597341371
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1597341371
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_44
timestamp 1597341371
transform 1 0 5152 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_32
timestamp 1597341371
transform 1 0 4048 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1597341371
transform 1 0 3588 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1597341371
transform 1 0 3956 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_63
timestamp 1597341371
transform 1 0 6900 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_56
timestamp 1597341371
transform 1 0 6256 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1597341371
transform 1 0 6808 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1597341371
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_87
timestamp 1597341371
transform 1 0 9108 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_75
timestamp 1597341371
transform 1 0 8004 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1597341371
transform 1 0 9660 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_118
timestamp 1597341371
transform 1 0 11960 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_106
timestamp 1597341371
transform 1 0 10856 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1597341371
transform 1 0 12512 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1597341371
transform 1 0 14812 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1597341371
transform 1 0 13708 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1597341371
transform 1 0 12604 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_168
timestamp 1597341371
transform 1 0 16560 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_156
timestamp 1597341371
transform 1 0 15456 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1597341371
transform 1 0 15364 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_187
timestamp 1597341371
transform 1 0 18308 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_180
timestamp 1597341371
transform 1 0 17664 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1597341371
transform 1 0 18216 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_218
timestamp 1597341371
transform 1 0 21160 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_211
timestamp 1597341371
transform 1 0 20516 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_199
timestamp 1597341371
transform 1 0 19412 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1597341371
transform 1 0 21068 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_242
timestamp 1597341371
transform 1 0 23368 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_230
timestamp 1597341371
transform 1 0 22264 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1597341371
transform 1 0 23920 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1597341371
transform 1 0 26220 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1597341371
transform 1 0 25116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1597341371
transform 1 0 24012 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_292
timestamp 1597341371
transform 1 0 27968 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_280
timestamp 1597341371
transform 1 0 26864 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1597341371
transform 1 0 26772 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1597341371
transform -1 0 28336 0 1 28832
box -38 -48 314 592
<< labels >>
rlabel metal2 s 18510 0 18566 800 6 CSB
port 0 nsew default input
rlabel metal2 s 24858 30871 24914 31671 6 RST
port 1 nsew default input
rlabel metal2 s 9218 0 9274 800 6 SCK
port 2 nsew default input
rlabel metal2 s 18 0 74 800 6 SDI
port 3 nsew default input
rlabel metal3 s 28727 24624 29527 24744 6 mask_rev_in[0]
port 4 nsew default input
rlabel metal3 s 0 27344 800 27464 6 mask_rev_in[1]
port 5 nsew default input
rlabel metal2 s 6366 30871 6422 31671 6 mask_rev_in[2]
port 6 nsew default input
rlabel metal2 s 27710 0 27766 800 6 mask_rev_in[3]
port 7 nsew default input
rlabel metal3 s 28727 11024 29527 11144 6 out
port 8 nsew default tristate
rlabel metal3 s 0 13608 800 13728 6 select
port 9 nsew default input
rlabel metal2 s 15658 30871 15714 31671 6 trap
port 10 nsew default input
rlabel metal5 s 1104 2768 28336 3088 6 VPWR
port 11 nsew default input
rlabel metal5 s 1104 4268 28336 4588 6 VGND
port 12 nsew default input
<< properties >>
string FIXED_BBOX 0 0 29527 31671
<< end >>

VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   # BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO AMUX2_3V
   CLASS BLOCK ;
   FOREIGN AMUX2_3V ;
   ORIGIN -0.5000 -2.1000 ;
   SIZE 9.0000 BY 5.4000 ;
   PIN select
      PORT
         LAYER metal1 ;
	    RECT 3.3000 4.0000 4.1000 4.4000 ;
      END
   END select
   PIN VDD
      PORT
         LAYER metal1 ;
	    RECT 0.5000 2.5000 0.9000 7.5000 ;
	    RECT 3.6000 2.5000 4.0000 3.6000 ;
	    RECT 0.5000 2.2000 4.0000 2.5000 ;
	    RECT 0.5000 2.1000 0.9000 2.2000 ;
      END
   END VDD
   PIN I0
      PORT
         LAYER metal1 ;
	    RECT 1.7000 3.3000 2.1000 5.8000 ;
      END
   END I0
   PIN I1
      PORT
         LAYER metal1 ;
	    RECT 7.9000 3.3000 8.3000 5.8000 ;
      END
   END I1
   PIN VSS
      PORT
         LAYER metal1 ;
	    RECT 3.6000 6.5000 5.8000 6.8000 ;
	    RECT 3.6000 5.5000 4.0000 6.5000 ;
	    RECT 5.5000 2.5000 5.8000 6.5000 ;
	    RECT 9.1000 2.5000 9.5000 7.5000 ;
	    RECT 5.5000 2.2000 9.5000 2.5000 ;
	    RECT 9.1000 2.1000 9.5000 2.2000 ;
      END
   END VSS
   PIN out
      PORT
         LAYER metal1 ;
	    RECT 2.5000 7.1000 7.5000 7.5000 ;
	    RECT 2.5000 3.3000 2.9000 7.1000 ;
	    RECT 7.1000 3.3000 7.5000 7.1000 ;
      END
   END out
   OBS
         LAYER metal1 ;
	    RECT 4.4000 5.1000 4.8000 5.8000 ;
	    RECT 3.4000 4.7000 5.0000 5.1000 ;
	    RECT 4.4000 3.3000 4.8000 4.7000 ;
   END
END AMUX2_3V

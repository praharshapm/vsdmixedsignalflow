VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AMUX2_3V
  CLASS CORE ;
  FOREIGN AMUX2_3V ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.060 BY 5.440 ;
  SITE unithddbl ;
  PIN select
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.644000 ;
    PORT
      LAYER li1 ;
        RECT 2.820 1.910 3.620 2.310 ;
    END
  END select
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 0.400 0.400 5.440 ;
        RECT 3.120 0.400 3.520 1.510 ;
        RECT 0.000 0.100 3.520 0.400 ;
        RECT 0.000 0.000 0.400 0.100 ;
    END
  END VDD
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.143100 ;
    PORT
      LAYER li1 ;
        RECT 1.200 1.200 1.610 3.720 ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.143100 ;
    PORT
      LAYER li1 ;
        RECT 7.450 1.200 7.850 3.720 ;
    END
  END I1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 3.120 4.430 5.330 4.730 ;
        RECT 3.120 3.420 3.520 4.430 ;
        RECT 5.030 0.400 5.330 4.430 ;
        RECT 8.660 0.400 9.060 5.440 ;
        RECT 5.030 0.100 9.060 0.400 ;
        RECT 8.660 0.000 9.060 0.100 ;
    END
  END VSS
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.270100 ;
    PORT
      LAYER li1 ;
        RECT 2.010 5.030 7.050 5.440 ;
        RECT 2.010 1.200 2.410 5.030 ;
        RECT 6.640 1.200 7.050 5.030 ;
    END
  END out
  OBS
      LAYER li1 ;
        RECT 3.920 3.020 4.330 3.720 ;
        RECT 2.920 2.610 4.530 3.020 ;
        RECT 3.920 1.200 4.330 2.610 ;
  END
END AMUX2_3V
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AMUX2_3V
  CLASS CORE ;
  FOREIGN AMUX2_3V ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 5.440 ;
  SITE unithddbl ;
  PIN select
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.648000 ;
    PORT
      LAYER li1 ;
        RECT 2.450 2.450 2.800 2.720 ;
    END
  END select
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.263600 ;
    PORT
      LAYER li1 ;
        RECT 6.890 3.620 7.610 4.400 ;
        RECT 6.940 2.260 7.340 3.620 ;
        RECT 6.890 1.500 7.610 2.260 ;
    END
  END I0
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.268000 ;
    PORT
      LAYER li1 ;
        RECT 1.130 3.620 1.850 4.400 ;
        RECT 6.040 3.620 6.610 4.400 ;
        RECT 1.210 2.280 1.600 3.620 ;
        RECT 1.130 1.500 1.850 2.280 ;
        RECT 6.160 2.260 6.560 3.620 ;
        RECT 6.040 1.500 6.610 2.260 ;
        RECT 1.200 1.190 1.600 1.500 ;
        RECT 6.160 1.190 6.560 1.500 ;
        RECT 1.200 1.020 6.560 1.190 ;
    END
  END out
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.036800 ;
    PORT
      LAYER li1 ;
        RECT 0.280 3.620 0.850 4.400 ;
        RECT 0.400 2.280 0.800 3.620 ;
        RECT 0.280 1.500 0.850 2.280 ;
    END
  END I1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.770 2.590 2.280 2.770 ;
        RECT 3.670 2.590 5.990 2.770 ;
        RECT 7.510 2.590 8.740 2.770 ;
        RECT 2.110 2.260 2.280 2.310 ;
        RECT 2.110 2.250 2.740 2.260 ;
        RECT 2.030 2.000 2.740 2.250 ;
        RECT 2.170 1.500 2.740 2.000 ;
      LAYER mcon ;
        RECT 1.910 2.590 2.090 2.770 ;
        RECT 3.820 2.590 4.000 2.770 ;
        RECT 4.310 2.590 4.490 2.770 ;
        RECT 4.800 2.590 4.980 2.770 ;
        RECT 5.290 2.590 5.470 2.770 ;
        RECT 5.780 2.590 5.960 2.770 ;
        RECT 7.660 2.590 7.840 2.770 ;
        RECT 8.150 2.590 8.330 2.770 ;
        RECT 2.110 2.140 2.280 2.310 ;
      LAYER met1 ;
        RECT 0.000 2.440 8.740 2.920 ;
        RECT 2.030 2.250 2.420 2.440 ;
        RECT 2.030 2.000 2.450 2.250 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.090 8.720 0.090 ;
      LAYER mcon ;
        RECT 0.150 -0.090 0.330 0.090 ;
        RECT 0.640 -0.090 0.820 0.090 ;
        RECT 1.130 -0.090 1.310 0.090 ;
        RECT 1.620 -0.090 1.800 0.090 ;
        RECT 2.110 -0.090 2.290 0.090 ;
        RECT 2.600 -0.090 2.780 0.090 ;
        RECT 3.090 -0.090 3.270 0.090 ;
        RECT 3.580 -0.090 3.760 0.090 ;
        RECT 4.070 -0.090 4.250 0.090 ;
        RECT 4.560 -0.090 4.740 0.090 ;
        RECT 5.050 -0.090 5.230 0.090 ;
        RECT 5.540 -0.090 5.720 0.090 ;
        RECT 6.030 -0.090 6.210 0.090 ;
        RECT 6.520 -0.090 6.700 0.090 ;
        RECT 7.010 -0.090 7.190 0.090 ;
        RECT 7.500 -0.090 7.680 0.090 ;
        RECT 7.990 -0.090 8.170 0.090 ;
        RECT 8.480 -0.090 8.660 0.090 ;
      LAYER met1 ;
        RECT 0.000 -0.240 8.720 0.240 ;
    END
  END VDD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000 5.350 8.740 5.530 ;
        RECT 2.290 4.400 2.690 5.350 ;
        RECT 2.170 3.620 2.740 4.400 ;
      LAYER mcon ;
        RECT 0.150 5.350 0.330 5.530 ;
        RECT 0.640 5.350 0.820 5.530 ;
        RECT 1.130 5.350 1.310 5.530 ;
        RECT 1.620 5.350 1.800 5.530 ;
        RECT 2.110 5.350 2.290 5.530 ;
        RECT 2.600 5.350 2.780 5.530 ;
        RECT 3.090 5.350 3.270 5.530 ;
        RECT 3.580 5.350 3.760 5.530 ;
        RECT 4.070 5.350 4.250 5.530 ;
        RECT 4.560 5.350 4.740 5.530 ;
        RECT 5.050 5.350 5.230 5.530 ;
        RECT 5.540 5.350 5.720 5.530 ;
        RECT 6.030 5.350 6.210 5.530 ;
        RECT 6.520 5.350 6.700 5.530 ;
        RECT 7.010 5.350 7.190 5.530 ;
        RECT 7.500 5.350 7.680 5.530 ;
        RECT 7.990 5.350 8.170 5.530 ;
        RECT 8.480 5.350 8.660 5.530 ;
      LAYER met1 ;
        RECT 0.000 5.200 8.740 5.680 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT 3.020 3.620 3.740 4.400 ;
        RECT 3.100 3.450 3.500 3.620 ;
        RECT 2.470 3.440 3.500 3.450 ;
        RECT 2.470 3.300 3.600 3.440 ;
        RECT 2.220 3.080 3.600 3.300 ;
        RECT 2.220 3.050 3.500 3.080 ;
        RECT 2.220 2.940 2.570 3.050 ;
        RECT 2.920 3.040 3.500 3.050 ;
        RECT 3.100 2.260 3.500 3.040 ;
        RECT 3.020 1.500 3.740 2.260 ;
  END
END AMUX2_3V
END LIBRARY


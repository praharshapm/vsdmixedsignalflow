magic
tech sky130A
magscale 1 2
timestamp 1598931070
<< locali >>
rect 18521 7735 18555 7837
rect 13553 7191 13587 7497
rect 14013 4539 14047 4641
<< viali >>
rect 23673 27421 23707 27455
rect 23029 27353 23063 27387
rect 23121 27081 23155 27115
rect 14105 16541 14139 16575
rect 15669 16541 15703 16575
rect 15485 16473 15519 16507
rect 16037 16473 16071 16507
rect 14289 16405 14323 16439
rect 14197 15997 14231 16031
rect 14473 15997 14507 16031
rect 16221 15997 16255 16031
rect 16497 15929 16531 15963
rect 13921 15861 13955 15895
rect 16865 15861 16899 15895
rect 17325 15861 17359 15895
rect 13921 15657 13955 15691
rect 16773 15521 16807 15555
rect 12725 15453 12759 15487
rect 15669 15453 15703 15487
rect 17233 15453 17267 15487
rect 17417 15453 17451 15487
rect 17785 15453 17819 15487
rect 17969 15453 18003 15487
rect 19441 15453 19475 15487
rect 15485 15385 15519 15419
rect 16037 15385 16071 15419
rect 12909 15317 12943 15351
rect 13277 15317 13311 15351
rect 14197 15317 14231 15351
rect 14657 15317 14691 15351
rect 16405 15317 16439 15351
rect 18521 15317 18555 15351
rect 19073 15317 19107 15351
rect 12817 15113 12851 15147
rect 15393 15113 15427 15147
rect 16313 15113 16347 15147
rect 14657 15045 14691 15079
rect 17141 15045 17175 15079
rect 18521 15045 18555 15079
rect 18797 15045 18831 15079
rect 13829 14977 13863 15011
rect 14289 14977 14323 15011
rect 15577 14977 15611 15011
rect 16589 14977 16623 15011
rect 16681 14977 16715 15011
rect 19441 14977 19475 15011
rect 20361 14909 20395 14943
rect 20637 14909 20671 14943
rect 22385 14909 22419 14943
rect 13645 14773 13679 14807
rect 17509 14773 17543 14807
rect 19901 14773 19935 14807
rect 14565 14569 14599 14603
rect 14933 14569 14967 14603
rect 17417 14569 17451 14603
rect 21373 14569 21407 14603
rect 21649 14569 21683 14603
rect 16497 14501 16531 14535
rect 17141 14501 17175 14535
rect 11897 14433 11931 14467
rect 15853 14365 15887 14399
rect 16221 14365 16255 14399
rect 16497 14365 16531 14399
rect 18245 14365 18279 14399
rect 18613 14365 18647 14399
rect 18797 14365 18831 14399
rect 19257 14365 19291 14399
rect 19349 14365 19383 14399
rect 21189 14365 21223 14399
rect 12173 14297 12207 14331
rect 13921 14297 13955 14331
rect 19901 14297 19935 14331
rect 17969 14229 18003 14263
rect 20361 14229 20395 14263
rect 11621 14025 11655 14059
rect 14565 14025 14599 14059
rect 17693 14025 17727 14059
rect 19901 14025 19935 14059
rect 20913 14025 20947 14059
rect 11897 13957 11931 13991
rect 12633 13957 12667 13991
rect 16405 13957 16439 13991
rect 18429 13957 18463 13991
rect 8585 13889 8619 13923
rect 13093 13889 13127 13923
rect 13277 13889 13311 13923
rect 13461 13889 13495 13923
rect 14105 13889 14139 13923
rect 14841 13889 14875 13923
rect 15117 13889 15151 13923
rect 16681 13889 16715 13923
rect 19073 13889 19107 13923
rect 19441 13889 19475 13923
rect 20453 13889 20487 13923
rect 13921 13821 13955 13855
rect 15577 13821 15611 13855
rect 18889 13821 18923 13855
rect 19349 13821 19383 13855
rect 8769 13753 8803 13787
rect 14933 13753 14967 13787
rect 20637 13753 20671 13787
rect 11253 13685 11287 13719
rect 15853 13685 15887 13719
rect 21373 13685 21407 13719
rect 11989 13481 12023 13515
rect 14841 13481 14875 13515
rect 17325 13481 17359 13515
rect 20453 13481 20487 13515
rect 10885 13413 10919 13447
rect 14565 13413 14599 13447
rect 15761 13413 15795 13447
rect 16865 13413 16899 13447
rect 11621 13345 11655 13379
rect 12909 13345 12943 13379
rect 13829 13345 13863 13379
rect 15632 13345 15666 13379
rect 15853 13345 15887 13379
rect 16589 13345 16623 13379
rect 18889 13345 18923 13379
rect 20085 13345 20119 13379
rect 11253 13277 11287 13311
rect 13369 13277 13403 13311
rect 13737 13277 13771 13311
rect 17049 13277 17083 13311
rect 17141 13277 17175 13311
rect 19073 13277 19107 13311
rect 19257 13277 19291 13311
rect 19625 13277 19659 13311
rect 19717 13277 19751 13311
rect 22293 13277 22327 13311
rect 15485 13209 15519 13243
rect 16221 13209 16255 13243
rect 22569 13209 22603 13243
rect 24317 13209 24351 13243
rect 8585 13141 8619 13175
rect 12541 13141 12575 13175
rect 17969 13141 18003 13175
rect 18245 13141 18279 13175
rect 21097 13141 21131 13175
rect 21833 13141 21867 13175
rect 11253 12937 11287 12971
rect 11713 12937 11747 12971
rect 16221 12937 16255 12971
rect 16589 12937 16623 12971
rect 16957 12937 16991 12971
rect 19257 12937 19291 12971
rect 20913 12937 20947 12971
rect 21465 12937 21499 12971
rect 23949 12937 23983 12971
rect 14197 12869 14231 12903
rect 20177 12869 20211 12903
rect 23029 12869 23063 12903
rect 13277 12801 13311 12835
rect 13553 12801 13587 12835
rect 15301 12801 15335 12835
rect 15669 12801 15703 12835
rect 15853 12801 15887 12835
rect 18797 12801 18831 12835
rect 18889 12801 18923 12835
rect 19073 12801 19107 12835
rect 22201 12801 22235 12835
rect 22569 12801 22603 12835
rect 12081 12733 12115 12767
rect 12909 12733 12943 12767
rect 13829 12733 13863 12767
rect 15209 12733 15243 12767
rect 19809 12733 19843 12767
rect 22661 12733 22695 12767
rect 18521 12665 18555 12699
rect 22017 12665 22051 12699
rect 14749 12597 14783 12631
rect 17233 12597 17267 12631
rect 17693 12597 17727 12631
rect 20637 12597 20671 12631
rect 13369 12393 13403 12427
rect 17049 12393 17083 12427
rect 19625 12393 19659 12427
rect 20177 12393 20211 12427
rect 22569 12393 22603 12427
rect 15761 12325 15795 12359
rect 11069 12257 11103 12291
rect 18337 12257 18371 12291
rect 22201 12257 22235 12291
rect 22845 12257 22879 12291
rect 23949 12257 23983 12291
rect 14197 12189 14231 12223
rect 15485 12189 15519 12223
rect 16405 12189 16439 12223
rect 16497 12189 16531 12223
rect 17601 12189 17635 12223
rect 17785 12189 17819 12223
rect 18245 12189 18279 12223
rect 19349 12189 19383 12223
rect 19441 12189 19475 12223
rect 21741 12189 21775 12223
rect 21925 12189 21959 12223
rect 11345 12121 11379 12155
rect 13093 12121 13127 12155
rect 10701 12053 10735 12087
rect 13829 12053 13863 12087
rect 14657 12053 14691 12087
rect 18889 12053 18923 12087
rect 21097 12053 21131 12087
rect 23489 12053 23523 12087
rect 24317 11917 24351 11951
rect 10701 11849 10735 11883
rect 11161 11849 11195 11883
rect 11437 11849 11471 11883
rect 14473 11849 14507 11883
rect 17049 11849 17083 11883
rect 22569 11849 22603 11883
rect 11805 11781 11839 11815
rect 12633 11781 12667 11815
rect 22937 11781 22971 11815
rect 8125 11713 8159 11747
rect 13185 11713 13219 11747
rect 13277 11713 13311 11747
rect 13461 11713 13495 11747
rect 14105 11713 14139 11747
rect 15209 11713 15243 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 18705 11713 18739 11747
rect 18889 11713 18923 11747
rect 19349 11713 19383 11747
rect 19441 11713 19475 11747
rect 21741 11713 21775 11747
rect 8033 11645 8067 11679
rect 13921 11645 13955 11679
rect 14749 11645 14783 11679
rect 15853 11645 15887 11679
rect 16129 11645 16163 11679
rect 18429 11645 18463 11679
rect 20913 11645 20947 11679
rect 21465 11645 21499 11679
rect 21925 11645 21959 11679
rect 25053 11645 25087 11679
rect 19809 11577 19843 11611
rect 8309 11509 8343 11543
rect 16497 11509 16531 11543
rect 17509 11509 17543 11543
rect 20361 11509 20395 11543
rect 22293 11509 22327 11543
rect 11069 11305 11103 11339
rect 12909 11305 12943 11339
rect 13277 11305 13311 11339
rect 15945 11305 15979 11339
rect 18061 11305 18095 11339
rect 18429 11305 18463 11339
rect 19533 11305 19567 11339
rect 19901 11305 19935 11339
rect 12081 11237 12115 11271
rect 13737 11237 13771 11271
rect 14473 11237 14507 11271
rect 16773 11237 16807 11271
rect 18797 11237 18831 11271
rect 12449 11169 12483 11203
rect 14105 11169 14139 11203
rect 19625 11169 19659 11203
rect 21833 11169 21867 11203
rect 22109 11169 22143 11203
rect 22477 11169 22511 11203
rect 6745 11101 6779 11135
rect 8125 11101 8159 11135
rect 8769 11101 8803 11135
rect 10885 11101 10919 11135
rect 11897 11101 11931 11135
rect 15485 11101 15519 11135
rect 16957 11101 16991 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 19404 11101 19438 11135
rect 21741 11101 21775 11135
rect 22569 11101 22603 11135
rect 7757 11033 7791 11067
rect 14841 11033 14875 11067
rect 19257 11033 19291 11067
rect 6929 10965 6963 10999
rect 9045 10965 9079 10999
rect 11621 10965 11655 10999
rect 15669 10965 15703 10999
rect 20453 10965 20487 10999
rect 6469 10761 6503 10795
rect 11069 10761 11103 10795
rect 13093 10761 13127 10795
rect 13461 10761 13495 10795
rect 17693 10761 17727 10795
rect 19441 10761 19475 10795
rect 19717 10761 19751 10795
rect 21833 10761 21867 10795
rect 12633 10693 12667 10727
rect 16221 10693 16255 10727
rect 17325 10693 17359 10727
rect 18981 10693 19015 10727
rect 20269 10693 20303 10727
rect 8401 10625 8435 10659
rect 8953 10625 8987 10659
rect 9137 10625 9171 10659
rect 10517 10625 10551 10659
rect 16773 10625 16807 10659
rect 18889 10625 18923 10659
rect 20913 10625 20947 10659
rect 21281 10625 21315 10659
rect 8309 10557 8343 10591
rect 13829 10557 13863 10591
rect 14105 10557 14139 10591
rect 15853 10557 15887 10591
rect 20821 10557 20855 10591
rect 21373 10557 21407 10591
rect 9321 10489 9355 10523
rect 10701 10489 10735 10523
rect 22845 10489 22879 10523
rect 7021 10421 7055 10455
rect 7481 10421 7515 10455
rect 7849 10421 7883 10455
rect 9873 10421 9907 10455
rect 11989 10421 12023 10455
rect 16957 10421 16991 10455
rect 22201 10421 22235 10455
rect 22477 10421 22511 10455
rect 6377 10217 6411 10251
rect 6929 10217 6963 10251
rect 9045 10217 9079 10251
rect 13001 10217 13035 10251
rect 13461 10217 13495 10251
rect 13921 10217 13955 10251
rect 14657 10217 14691 10251
rect 17509 10217 17543 10251
rect 18061 10217 18095 10251
rect 18981 10217 19015 10251
rect 19717 10217 19751 10251
rect 21465 10217 21499 10251
rect 21097 10149 21131 10183
rect 10425 10081 10459 10115
rect 17141 10081 17175 10115
rect 19073 10081 19107 10115
rect 21833 10081 21867 10115
rect 23857 10081 23891 10115
rect 6193 10013 6227 10047
rect 7665 10013 7699 10047
rect 7941 10013 7975 10047
rect 8033 10013 8067 10047
rect 8309 10013 8343 10047
rect 8585 10013 8619 10047
rect 13737 10013 13771 10047
rect 15669 10013 15703 10047
rect 16405 10013 16439 10047
rect 16865 10013 16899 10047
rect 18429 10013 18463 10047
rect 18852 10013 18886 10047
rect 7205 9945 7239 9979
rect 10701 9945 10735 9979
rect 12449 9945 12483 9979
rect 15485 9945 15519 9979
rect 16037 9945 16071 9979
rect 16681 9945 16715 9979
rect 18705 9945 18739 9979
rect 22109 9945 22143 9979
rect 10149 9877 10183 9911
rect 14197 9877 14231 9911
rect 19349 9877 19383 9911
rect 20269 9877 20303 9911
rect 5733 9673 5767 9707
rect 9781 9673 9815 9707
rect 11805 9673 11839 9707
rect 14197 9673 14231 9707
rect 15393 9673 15427 9707
rect 21557 9673 21591 9707
rect 22017 9673 22051 9707
rect 22661 9673 22695 9707
rect 6101 9605 6135 9639
rect 6469 9605 6503 9639
rect 9413 9605 9447 9639
rect 15025 9605 15059 9639
rect 17693 9605 17727 9639
rect 20269 9605 20303 9639
rect 10517 9537 10551 9571
rect 10701 9537 10735 9571
rect 10977 9537 11011 9571
rect 13093 9537 13127 9571
rect 14381 9537 14415 9571
rect 15945 9537 15979 9571
rect 16497 9537 16531 9571
rect 16681 9537 16715 9571
rect 18889 9537 18923 9571
rect 19073 9537 19107 9571
rect 19257 9537 19291 9571
rect 20416 9537 20450 9571
rect 21833 9537 21867 9571
rect 23029 9537 23063 9571
rect 7021 9469 7055 9503
rect 7297 9469 7331 9503
rect 9045 9469 9079 9503
rect 10057 9469 10091 9503
rect 11161 9469 11195 9503
rect 11437 9469 11471 9503
rect 15853 9469 15887 9503
rect 20637 9469 20671 9503
rect 22293 9469 22327 9503
rect 18705 9401 18739 9435
rect 20545 9401 20579 9435
rect 13461 9333 13495 9367
rect 16957 9333 16991 9367
rect 19809 9333 19843 9367
rect 20913 9333 20947 9367
rect 7665 9129 7699 9163
rect 8493 9129 8527 9163
rect 9229 9129 9263 9163
rect 10701 9129 10735 9163
rect 11345 9129 11379 9163
rect 15853 9129 15887 9163
rect 16129 9129 16163 9163
rect 16589 9129 16623 9163
rect 19165 9129 19199 9163
rect 19901 9129 19935 9163
rect 22293 9129 22327 9163
rect 6561 9061 6595 9095
rect 7021 9061 7055 9095
rect 22753 9061 22787 9095
rect 7389 8993 7423 9027
rect 10425 8993 10459 9027
rect 11897 8993 11931 9027
rect 12725 8993 12759 9027
rect 13691 8993 13725 9027
rect 14933 8993 14967 9027
rect 17141 8993 17175 9027
rect 18889 8993 18923 9027
rect 21097 8993 21131 9027
rect 6837 8925 6871 8959
rect 8401 8925 8435 8959
rect 10057 8925 10091 8959
rect 11253 8925 11287 8959
rect 13553 8925 13587 8959
rect 13829 8925 13863 8959
rect 16865 8925 16899 8959
rect 19717 8925 19751 8959
rect 21281 8925 21315 8959
rect 21741 8925 21775 8959
rect 21833 8925 21867 8959
rect 8217 8857 8251 8891
rect 9873 8857 9907 8891
rect 11069 8857 11103 8891
rect 13001 8857 13035 8891
rect 23121 8857 23155 8891
rect 6193 8789 6227 8823
rect 14381 8789 14415 8823
rect 20269 8789 20303 8823
rect 6101 8585 6135 8619
rect 10517 8585 10551 8619
rect 11805 8585 11839 8619
rect 17233 8585 17267 8619
rect 17693 8585 17727 8619
rect 18429 8585 18463 8619
rect 19073 8585 19107 8619
rect 21189 8585 21223 8619
rect 21557 8585 21591 8619
rect 22661 8585 22695 8619
rect 7665 8517 7699 8551
rect 8033 8517 8067 8551
rect 8493 8517 8527 8551
rect 14933 8517 14967 8551
rect 15393 8517 15427 8551
rect 7205 8449 7239 8483
rect 9321 8449 9355 8483
rect 11437 8449 11471 8483
rect 15853 8449 15887 8483
rect 18245 8449 18279 8483
rect 19441 8449 19475 8483
rect 19533 8449 19567 8483
rect 19717 8449 19751 8483
rect 20085 8449 20119 8483
rect 20278 8449 20312 8483
rect 21925 8449 21959 8483
rect 7113 8381 7147 8415
rect 9045 8381 9079 8415
rect 9505 8381 9539 8415
rect 10793 8381 10827 8415
rect 12909 8381 12943 8415
rect 13185 8381 13219 8415
rect 20637 8381 20671 8415
rect 10057 8313 10091 8347
rect 16957 8313 16991 8347
rect 6377 8245 6411 8279
rect 16221 8245 16255 8279
rect 22293 8245 22327 8279
rect 7113 8041 7147 8075
rect 9045 8041 9079 8075
rect 11253 8041 11287 8075
rect 13001 8041 13035 8075
rect 14197 8041 14231 8075
rect 15853 8041 15887 8075
rect 16221 8041 16255 8075
rect 17877 8041 17911 8075
rect 21373 8041 21407 8075
rect 10977 7973 11011 8007
rect 18337 7973 18371 8007
rect 19717 7973 19751 8007
rect 6837 7905 6871 7939
rect 8309 7905 8343 7939
rect 13829 7905 13863 7939
rect 18705 7905 18739 7939
rect 21557 7905 21591 7939
rect 22017 7905 22051 7939
rect 6469 7837 6503 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 9873 7837 9907 7871
rect 9965 7837 9999 7871
rect 10149 7837 10183 7871
rect 12541 7837 12575 7871
rect 13369 7837 13403 7871
rect 16681 7837 16715 7871
rect 18153 7837 18187 7871
rect 18521 7837 18555 7871
rect 18981 7837 19015 7871
rect 20453 7837 20487 7871
rect 21741 7837 21775 7871
rect 22109 7837 22143 7871
rect 7757 7769 7791 7803
rect 10609 7769 10643 7803
rect 17325 7769 17359 7803
rect 11621 7701 11655 7735
rect 12265 7701 12299 7735
rect 13553 7701 13587 7735
rect 18521 7701 18555 7735
rect 19349 7701 19383 7735
rect 20085 7701 20119 7735
rect 7021 7497 7055 7531
rect 7389 7497 7423 7531
rect 7849 7497 7883 7531
rect 10057 7497 10091 7531
rect 11621 7497 11655 7531
rect 13553 7497 13587 7531
rect 13645 7497 13679 7531
rect 16681 7497 16715 7531
rect 17325 7497 17359 7531
rect 17693 7497 17727 7531
rect 18245 7497 18279 7531
rect 20453 7497 20487 7531
rect 20821 7497 20855 7531
rect 22201 7497 22235 7531
rect 8493 7429 8527 7463
rect 9689 7429 9723 7463
rect 11253 7429 11287 7463
rect 12633 7429 12667 7463
rect 9137 7361 9171 7395
rect 10425 7361 10459 7395
rect 13277 7361 13311 7395
rect 21189 7429 21223 7463
rect 14749 7361 14783 7395
rect 14841 7361 14875 7395
rect 15209 7361 15243 7395
rect 15301 7361 15335 7395
rect 19073 7361 19107 7395
rect 19441 7361 19475 7395
rect 21833 7361 21867 7395
rect 19349 7293 19383 7327
rect 19901 7293 19935 7327
rect 8217 7157 8251 7191
rect 10609 7157 10643 7191
rect 10977 7157 11011 7191
rect 12081 7157 12115 7191
rect 13553 7157 13587 7191
rect 14197 7157 14231 7191
rect 15761 7157 15795 7191
rect 18705 7157 18739 7191
rect 8401 6953 8435 6987
rect 9321 6953 9355 6987
rect 10149 6953 10183 6987
rect 10885 6953 10919 6987
rect 13737 6953 13771 6987
rect 14565 6953 14599 6987
rect 16313 6953 16347 6987
rect 16865 6953 16899 6987
rect 17877 6953 17911 6987
rect 21189 6953 21223 6987
rect 8769 6885 8803 6919
rect 14289 6885 14323 6919
rect 11437 6817 11471 6851
rect 13461 6817 13495 6851
rect 15485 6817 15519 6851
rect 19993 6817 20027 6851
rect 6285 6749 6319 6783
rect 7481 6749 7515 6783
rect 7665 6749 7699 6783
rect 8033 6749 8067 6783
rect 10057 6749 10091 6783
rect 15577 6749 15611 6783
rect 16681 6749 16715 6783
rect 17693 6749 17727 6783
rect 18153 6749 18187 6783
rect 18613 6749 18647 6783
rect 19901 6749 19935 6783
rect 21465 6749 21499 6783
rect 21925 6749 21959 6783
rect 7021 6681 7055 6715
rect 11713 6681 11747 6715
rect 16037 6681 16071 6715
rect 6469 6613 6503 6647
rect 18889 6613 18923 6647
rect 20269 6613 20303 6647
rect 21649 6613 21683 6647
rect 22293 6613 22327 6647
rect 7205 6409 7239 6443
rect 9505 6409 9539 6443
rect 10701 6409 10735 6443
rect 14105 6409 14139 6443
rect 5365 6341 5399 6375
rect 5917 6341 5951 6375
rect 9781 6341 9815 6375
rect 11069 6341 11103 6375
rect 12633 6341 12667 6375
rect 15301 6341 15335 6375
rect 15669 6341 15703 6375
rect 16129 6341 16163 6375
rect 18337 6341 18371 6375
rect 5549 6273 5583 6307
rect 6285 6273 6319 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8769 6273 8803 6307
rect 9965 6273 9999 6307
rect 11345 6273 11379 6307
rect 11805 6273 11839 6307
rect 13093 6273 13127 6307
rect 13461 6273 13495 6307
rect 14381 6273 14415 6307
rect 14473 6273 14507 6307
rect 16957 6273 16991 6307
rect 19349 6273 19383 6307
rect 19717 6273 19751 6307
rect 7481 6205 7515 6239
rect 8861 6205 8895 6239
rect 10241 6205 10275 6239
rect 13553 6205 13587 6239
rect 16681 6205 16715 6239
rect 17141 6205 17175 6239
rect 19441 6205 19475 6239
rect 19625 6205 19659 6239
rect 20177 6205 20211 6239
rect 20729 6205 20763 6239
rect 21005 6205 21039 6239
rect 22753 6205 22787 6239
rect 11529 6137 11563 6171
rect 14657 6069 14691 6103
rect 17417 6069 17451 6103
rect 18981 6069 19015 6103
rect 5365 5865 5399 5899
rect 5825 5865 5859 5899
rect 9045 5865 9079 5899
rect 10977 5865 11011 5899
rect 14381 5865 14415 5899
rect 18521 5865 18555 5899
rect 20545 5865 20579 5899
rect 10609 5797 10643 5831
rect 17969 5797 18003 5831
rect 6745 5729 6779 5763
rect 7021 5729 7055 5763
rect 8769 5729 8803 5763
rect 11989 5729 12023 5763
rect 13645 5729 13679 5763
rect 16037 5729 16071 5763
rect 16589 5729 16623 5763
rect 18797 5729 18831 5763
rect 20177 5729 20211 5763
rect 21097 5729 21131 5763
rect 21833 5729 21867 5763
rect 22017 5729 22051 5763
rect 9965 5661 9999 5695
rect 12817 5661 12851 5695
rect 12909 5661 12943 5695
rect 14197 5661 14231 5695
rect 16129 5661 16163 5695
rect 16497 5661 16531 5695
rect 17417 5661 17451 5695
rect 17785 5661 17819 5695
rect 18889 5661 18923 5695
rect 19625 5661 19659 5695
rect 21741 5661 21775 5695
rect 22109 5661 22143 5695
rect 11253 5593 11287 5627
rect 11437 5593 11471 5627
rect 11621 5593 11655 5627
rect 13369 5593 13403 5627
rect 15485 5593 15519 5627
rect 19349 5593 19383 5627
rect 6469 5525 6503 5559
rect 11529 5525 11563 5559
rect 12541 5525 12575 5559
rect 14657 5525 14691 5559
rect 16957 5525 16991 5559
rect 6469 5321 6503 5355
rect 7389 5321 7423 5355
rect 8125 5321 8159 5355
rect 14289 5321 14323 5355
rect 17325 5321 17359 5355
rect 18337 5321 18371 5355
rect 21097 5321 21131 5355
rect 21833 5321 21867 5355
rect 7849 5253 7883 5287
rect 8677 5253 8711 5287
rect 11621 5253 11655 5287
rect 16681 5253 16715 5287
rect 18981 5253 19015 5287
rect 21373 5253 21407 5287
rect 7021 5185 7055 5219
rect 9505 5185 9539 5219
rect 9689 5185 9723 5219
rect 11161 5185 11195 5219
rect 11253 5185 11287 5219
rect 12633 5185 12667 5219
rect 12909 5185 12943 5219
rect 13369 5185 13403 5219
rect 14657 5185 14691 5219
rect 15301 5185 15335 5219
rect 15669 5185 15703 5219
rect 16241 5185 16275 5219
rect 16957 5185 16991 5219
rect 9229 5117 9263 5151
rect 12725 5117 12759 5151
rect 16129 5117 16163 5151
rect 18705 5117 18739 5151
rect 20729 5117 20763 5151
rect 11897 5049 11931 5083
rect 10241 4981 10275 5015
rect 13921 4981 13955 5015
rect 6837 4777 6871 4811
rect 7573 4777 7607 4811
rect 9137 4777 9171 4811
rect 11897 4777 11931 4811
rect 13921 4777 13955 4811
rect 14657 4777 14691 4811
rect 18337 4777 18371 4811
rect 19809 4777 19843 4811
rect 20177 4777 20211 4811
rect 21557 4777 21591 4811
rect 18797 4709 18831 4743
rect 19165 4709 19199 4743
rect 21189 4709 21223 4743
rect 7941 4641 7975 4675
rect 10057 4641 10091 4675
rect 14013 4641 14047 4675
rect 16037 4641 16071 4675
rect 17785 4641 17819 4675
rect 8361 4573 8395 4607
rect 10333 4573 10367 4607
rect 10793 4573 10827 4607
rect 10977 4573 11011 4607
rect 11345 4573 11379 4607
rect 11529 4573 11563 4607
rect 13001 4573 13035 4607
rect 14206 4573 14240 4607
rect 15761 4573 15795 4607
rect 18613 4573 18647 4607
rect 19625 4573 19659 4607
rect 8217 4505 8251 4539
rect 13093 4505 13127 4539
rect 13553 4505 13587 4539
rect 14013 4505 14047 4539
rect 7113 4437 7147 4471
rect 8493 4437 8527 4471
rect 14381 4437 14415 4471
rect 20453 4437 20487 4471
rect 10701 4233 10735 4267
rect 11989 4233 12023 4267
rect 14933 4233 14967 4267
rect 15485 4233 15519 4267
rect 18705 4233 18739 4267
rect 19349 4233 19383 4267
rect 11621 4165 11655 4199
rect 12725 4165 12759 4199
rect 14289 4165 14323 4199
rect 7665 4097 7699 4131
rect 8309 4097 8343 4131
rect 12817 4097 12851 4131
rect 14013 4097 14047 4131
rect 16773 4097 16807 4131
rect 18245 4097 18279 4131
rect 18521 4097 18555 4131
rect 19625 4097 19659 4131
rect 20085 4097 20119 4131
rect 8585 4029 8619 4063
rect 10333 4029 10367 4063
rect 11345 4029 11379 4063
rect 14657 4029 14691 4063
rect 17601 4029 17635 4063
rect 14454 3961 14488 3995
rect 16589 3961 16623 3995
rect 17233 3961 17267 3995
rect 18337 3961 18371 3995
rect 6469 3893 6503 3927
rect 7205 3893 7239 3927
rect 8033 3893 8067 3927
rect 14565 3893 14599 3927
rect 15761 3893 15795 3927
rect 19809 3893 19843 3927
rect 20453 3893 20487 3927
rect 7021 3689 7055 3723
rect 11805 3689 11839 3723
rect 14657 3689 14691 3723
rect 18153 3689 18187 3723
rect 20085 3689 20119 3723
rect 14381 3621 14415 3655
rect 19165 3621 19199 3655
rect 7757 3553 7791 3587
rect 8677 3553 8711 3587
rect 10149 3553 10183 3587
rect 10977 3553 11011 3587
rect 11437 3553 11471 3587
rect 17509 3553 17543 3587
rect 8585 3485 8619 3519
rect 11253 3485 11287 3519
rect 12541 3485 12575 3519
rect 13093 3485 13127 3519
rect 13553 3485 13587 3519
rect 15761 3485 15795 3519
rect 16129 3485 16163 3519
rect 18705 3485 18739 3519
rect 7849 3417 7883 3451
rect 10425 3417 10459 3451
rect 12173 3417 12207 3451
rect 7389 3349 7423 3383
rect 9137 3349 9171 3383
rect 12633 3349 12667 3383
rect 14013 3349 14047 3383
rect 18889 3349 18923 3383
rect 19625 3349 19659 3383
rect 6469 3145 6503 3179
rect 7481 3145 7515 3179
rect 7849 3145 7883 3179
rect 8401 3145 8435 3179
rect 8769 3145 8803 3179
rect 15485 3145 15519 3179
rect 19165 3145 19199 3179
rect 19533 3145 19567 3179
rect 9781 3077 9815 3111
rect 11529 3077 11563 3111
rect 13185 3077 13219 3111
rect 14933 3077 14967 3111
rect 16405 3077 16439 3111
rect 18705 3077 18739 3111
rect 7297 3009 7331 3043
rect 9137 3009 9171 3043
rect 16957 3009 16991 3043
rect 18245 3009 18279 3043
rect 9505 2941 9539 2975
rect 12909 2941 12943 2975
rect 15761 2941 15795 2975
rect 18429 2873 18463 2907
rect 12081 2805 12115 2839
rect 17509 2805 17543 2839
rect 7665 2601 7699 2635
rect 9045 2601 9079 2635
rect 10149 2601 10183 2635
rect 10517 2601 10551 2635
rect 11437 2601 11471 2635
rect 12909 2601 12943 2635
rect 13277 2601 13311 2635
rect 17049 2601 17083 2635
rect 18889 2601 18923 2635
rect 8677 2533 8711 2567
rect 12265 2533 12299 2567
rect 13921 2533 13955 2567
rect 17417 2533 17451 2567
rect 17969 2533 18003 2567
rect 10885 2465 10919 2499
rect 7389 2397 7423 2431
rect 8309 2397 8343 2431
rect 9965 2397 9999 2431
rect 11161 2397 11195 2431
rect 11253 2397 11287 2431
rect 13829 2397 13863 2431
rect 14105 2397 14139 2431
rect 15117 2397 15151 2431
rect 16313 2397 16347 2431
rect 18705 2397 18739 2431
rect 19165 2397 19199 2431
rect 15669 2329 15703 2363
rect 16773 2329 16807 2363
rect 9321 2261 9355 2295
rect 14289 2261 14323 2295
<< metal1 >>
rect 1104 29402 28336 29424
rect 1104 29350 1782 29402
rect 1834 29350 1846 29402
rect 1898 29350 1910 29402
rect 1962 29350 1974 29402
rect 2026 29350 4782 29402
rect 4834 29350 4846 29402
rect 4898 29350 4910 29402
rect 4962 29350 4974 29402
rect 5026 29350 7782 29402
rect 7834 29350 7846 29402
rect 7898 29350 7910 29402
rect 7962 29350 7974 29402
rect 8026 29350 10782 29402
rect 10834 29350 10846 29402
rect 10898 29350 10910 29402
rect 10962 29350 10974 29402
rect 11026 29350 13782 29402
rect 13834 29350 13846 29402
rect 13898 29350 13910 29402
rect 13962 29350 13974 29402
rect 14026 29350 16782 29402
rect 16834 29350 16846 29402
rect 16898 29350 16910 29402
rect 16962 29350 16974 29402
rect 17026 29350 19782 29402
rect 19834 29350 19846 29402
rect 19898 29350 19910 29402
rect 19962 29350 19974 29402
rect 20026 29350 22782 29402
rect 22834 29350 22846 29402
rect 22898 29350 22910 29402
rect 22962 29350 22974 29402
rect 23026 29350 25782 29402
rect 25834 29350 25846 29402
rect 25898 29350 25910 29402
rect 25962 29350 25974 29402
rect 26026 29350 28336 29402
rect 1104 29328 28336 29350
rect 1104 28858 28336 28880
rect 1104 28806 3282 28858
rect 3334 28806 3346 28858
rect 3398 28806 3410 28858
rect 3462 28806 3474 28858
rect 3526 28806 6282 28858
rect 6334 28806 6346 28858
rect 6398 28806 6410 28858
rect 6462 28806 6474 28858
rect 6526 28806 9282 28858
rect 9334 28806 9346 28858
rect 9398 28806 9410 28858
rect 9462 28806 9474 28858
rect 9526 28806 12282 28858
rect 12334 28806 12346 28858
rect 12398 28806 12410 28858
rect 12462 28806 12474 28858
rect 12526 28806 15282 28858
rect 15334 28806 15346 28858
rect 15398 28806 15410 28858
rect 15462 28806 15474 28858
rect 15526 28806 18282 28858
rect 18334 28806 18346 28858
rect 18398 28806 18410 28858
rect 18462 28806 18474 28858
rect 18526 28806 21282 28858
rect 21334 28806 21346 28858
rect 21398 28806 21410 28858
rect 21462 28806 21474 28858
rect 21526 28806 24282 28858
rect 24334 28806 24346 28858
rect 24398 28806 24410 28858
rect 24462 28806 24474 28858
rect 24526 28806 27282 28858
rect 27334 28806 27346 28858
rect 27398 28806 27410 28858
rect 27462 28806 27474 28858
rect 27526 28806 28336 28858
rect 1104 28784 28336 28806
rect 1104 28314 28336 28336
rect 1104 28262 1782 28314
rect 1834 28262 1846 28314
rect 1898 28262 1910 28314
rect 1962 28262 1974 28314
rect 2026 28262 4782 28314
rect 4834 28262 4846 28314
rect 4898 28262 4910 28314
rect 4962 28262 4974 28314
rect 5026 28262 7782 28314
rect 7834 28262 7846 28314
rect 7898 28262 7910 28314
rect 7962 28262 7974 28314
rect 8026 28262 10782 28314
rect 10834 28262 10846 28314
rect 10898 28262 10910 28314
rect 10962 28262 10974 28314
rect 11026 28262 13782 28314
rect 13834 28262 13846 28314
rect 13898 28262 13910 28314
rect 13962 28262 13974 28314
rect 14026 28262 16782 28314
rect 16834 28262 16846 28314
rect 16898 28262 16910 28314
rect 16962 28262 16974 28314
rect 17026 28262 19782 28314
rect 19834 28262 19846 28314
rect 19898 28262 19910 28314
rect 19962 28262 19974 28314
rect 20026 28262 22782 28314
rect 22834 28262 22846 28314
rect 22898 28262 22910 28314
rect 22962 28262 22974 28314
rect 23026 28262 25782 28314
rect 25834 28262 25846 28314
rect 25898 28262 25910 28314
rect 25962 28262 25974 28314
rect 26026 28262 28336 28314
rect 1104 28240 28336 28262
rect 1104 27770 28336 27792
rect 1104 27718 3282 27770
rect 3334 27718 3346 27770
rect 3398 27718 3410 27770
rect 3462 27718 3474 27770
rect 3526 27718 6282 27770
rect 6334 27718 6346 27770
rect 6398 27718 6410 27770
rect 6462 27718 6474 27770
rect 6526 27718 9282 27770
rect 9334 27718 9346 27770
rect 9398 27718 9410 27770
rect 9462 27718 9474 27770
rect 9526 27718 12282 27770
rect 12334 27718 12346 27770
rect 12398 27718 12410 27770
rect 12462 27718 12474 27770
rect 12526 27718 15282 27770
rect 15334 27718 15346 27770
rect 15398 27718 15410 27770
rect 15462 27718 15474 27770
rect 15526 27718 18282 27770
rect 18334 27718 18346 27770
rect 18398 27718 18410 27770
rect 18462 27718 18474 27770
rect 18526 27718 21282 27770
rect 21334 27718 21346 27770
rect 21398 27718 21410 27770
rect 21462 27718 21474 27770
rect 21526 27718 24282 27770
rect 24334 27718 24346 27770
rect 24398 27718 24410 27770
rect 24462 27718 24474 27770
rect 24526 27718 27282 27770
rect 27334 27718 27346 27770
rect 27398 27718 27410 27770
rect 27462 27718 27474 27770
rect 27526 27718 28336 27770
rect 1104 27696 28336 27718
rect 23106 27412 23112 27464
rect 23164 27452 23170 27464
rect 23661 27455 23719 27461
rect 23661 27452 23673 27455
rect 23164 27424 23673 27452
rect 23164 27412 23170 27424
rect 23661 27421 23673 27424
rect 23707 27452 23719 27455
rect 24578 27452 24584 27464
rect 23707 27424 24584 27452
rect 23707 27421 23719 27424
rect 23661 27415 23719 27421
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 21634 27344 21640 27396
rect 21692 27384 21698 27396
rect 23017 27387 23075 27393
rect 23017 27384 23029 27387
rect 21692 27356 23029 27384
rect 21692 27344 21698 27356
rect 23017 27353 23029 27356
rect 23063 27353 23075 27387
rect 23017 27347 23075 27353
rect 1104 27226 28336 27248
rect 1104 27174 1782 27226
rect 1834 27174 1846 27226
rect 1898 27174 1910 27226
rect 1962 27174 1974 27226
rect 2026 27174 4782 27226
rect 4834 27174 4846 27226
rect 4898 27174 4910 27226
rect 4962 27174 4974 27226
rect 5026 27174 7782 27226
rect 7834 27174 7846 27226
rect 7898 27174 7910 27226
rect 7962 27174 7974 27226
rect 8026 27174 10782 27226
rect 10834 27174 10846 27226
rect 10898 27174 10910 27226
rect 10962 27174 10974 27226
rect 11026 27174 13782 27226
rect 13834 27174 13846 27226
rect 13898 27174 13910 27226
rect 13962 27174 13974 27226
rect 14026 27174 16782 27226
rect 16834 27174 16846 27226
rect 16898 27174 16910 27226
rect 16962 27174 16974 27226
rect 17026 27174 19782 27226
rect 19834 27174 19846 27226
rect 19898 27174 19910 27226
rect 19962 27174 19974 27226
rect 20026 27174 22782 27226
rect 22834 27174 22846 27226
rect 22898 27174 22910 27226
rect 22962 27174 22974 27226
rect 23026 27174 25782 27226
rect 25834 27174 25846 27226
rect 25898 27174 25910 27226
rect 25962 27174 25974 27226
rect 26026 27174 28336 27226
rect 1104 27152 28336 27174
rect 23106 27112 23112 27124
rect 23067 27084 23112 27112
rect 23106 27072 23112 27084
rect 23164 27072 23170 27124
rect 1104 26682 28336 26704
rect 1104 26630 3282 26682
rect 3334 26630 3346 26682
rect 3398 26630 3410 26682
rect 3462 26630 3474 26682
rect 3526 26630 6282 26682
rect 6334 26630 6346 26682
rect 6398 26630 6410 26682
rect 6462 26630 6474 26682
rect 6526 26630 9282 26682
rect 9334 26630 9346 26682
rect 9398 26630 9410 26682
rect 9462 26630 9474 26682
rect 9526 26630 12282 26682
rect 12334 26630 12346 26682
rect 12398 26630 12410 26682
rect 12462 26630 12474 26682
rect 12526 26630 15282 26682
rect 15334 26630 15346 26682
rect 15398 26630 15410 26682
rect 15462 26630 15474 26682
rect 15526 26630 18282 26682
rect 18334 26630 18346 26682
rect 18398 26630 18410 26682
rect 18462 26630 18474 26682
rect 18526 26630 21282 26682
rect 21334 26630 21346 26682
rect 21398 26630 21410 26682
rect 21462 26630 21474 26682
rect 21526 26630 24282 26682
rect 24334 26630 24346 26682
rect 24398 26630 24410 26682
rect 24462 26630 24474 26682
rect 24526 26630 27282 26682
rect 27334 26630 27346 26682
rect 27398 26630 27410 26682
rect 27462 26630 27474 26682
rect 27526 26630 28336 26682
rect 1104 26608 28336 26630
rect 1104 26138 28336 26160
rect 1104 26086 1782 26138
rect 1834 26086 1846 26138
rect 1898 26086 1910 26138
rect 1962 26086 1974 26138
rect 2026 26086 4782 26138
rect 4834 26086 4846 26138
rect 4898 26086 4910 26138
rect 4962 26086 4974 26138
rect 5026 26086 7782 26138
rect 7834 26086 7846 26138
rect 7898 26086 7910 26138
rect 7962 26086 7974 26138
rect 8026 26086 10782 26138
rect 10834 26086 10846 26138
rect 10898 26086 10910 26138
rect 10962 26086 10974 26138
rect 11026 26086 13782 26138
rect 13834 26086 13846 26138
rect 13898 26086 13910 26138
rect 13962 26086 13974 26138
rect 14026 26086 16782 26138
rect 16834 26086 16846 26138
rect 16898 26086 16910 26138
rect 16962 26086 16974 26138
rect 17026 26086 19782 26138
rect 19834 26086 19846 26138
rect 19898 26086 19910 26138
rect 19962 26086 19974 26138
rect 20026 26086 22782 26138
rect 22834 26086 22846 26138
rect 22898 26086 22910 26138
rect 22962 26086 22974 26138
rect 23026 26086 25782 26138
rect 25834 26086 25846 26138
rect 25898 26086 25910 26138
rect 25962 26086 25974 26138
rect 26026 26086 28336 26138
rect 1104 26064 28336 26086
rect 1104 25594 28336 25616
rect 1104 25542 3282 25594
rect 3334 25542 3346 25594
rect 3398 25542 3410 25594
rect 3462 25542 3474 25594
rect 3526 25542 6282 25594
rect 6334 25542 6346 25594
rect 6398 25542 6410 25594
rect 6462 25542 6474 25594
rect 6526 25542 9282 25594
rect 9334 25542 9346 25594
rect 9398 25542 9410 25594
rect 9462 25542 9474 25594
rect 9526 25542 12282 25594
rect 12334 25542 12346 25594
rect 12398 25542 12410 25594
rect 12462 25542 12474 25594
rect 12526 25542 15282 25594
rect 15334 25542 15346 25594
rect 15398 25542 15410 25594
rect 15462 25542 15474 25594
rect 15526 25542 18282 25594
rect 18334 25542 18346 25594
rect 18398 25542 18410 25594
rect 18462 25542 18474 25594
rect 18526 25542 21282 25594
rect 21334 25542 21346 25594
rect 21398 25542 21410 25594
rect 21462 25542 21474 25594
rect 21526 25542 24282 25594
rect 24334 25542 24346 25594
rect 24398 25542 24410 25594
rect 24462 25542 24474 25594
rect 24526 25542 27282 25594
rect 27334 25542 27346 25594
rect 27398 25542 27410 25594
rect 27462 25542 27474 25594
rect 27526 25542 28336 25594
rect 1104 25520 28336 25542
rect 1104 25050 28336 25072
rect 1104 24998 1782 25050
rect 1834 24998 1846 25050
rect 1898 24998 1910 25050
rect 1962 24998 1974 25050
rect 2026 24998 4782 25050
rect 4834 24998 4846 25050
rect 4898 24998 4910 25050
rect 4962 24998 4974 25050
rect 5026 24998 7782 25050
rect 7834 24998 7846 25050
rect 7898 24998 7910 25050
rect 7962 24998 7974 25050
rect 8026 24998 10782 25050
rect 10834 24998 10846 25050
rect 10898 24998 10910 25050
rect 10962 24998 10974 25050
rect 11026 24998 13782 25050
rect 13834 24998 13846 25050
rect 13898 24998 13910 25050
rect 13962 24998 13974 25050
rect 14026 24998 16782 25050
rect 16834 24998 16846 25050
rect 16898 24998 16910 25050
rect 16962 24998 16974 25050
rect 17026 24998 19782 25050
rect 19834 24998 19846 25050
rect 19898 24998 19910 25050
rect 19962 24998 19974 25050
rect 20026 24998 22782 25050
rect 22834 24998 22846 25050
rect 22898 24998 22910 25050
rect 22962 24998 22974 25050
rect 23026 24998 25782 25050
rect 25834 24998 25846 25050
rect 25898 24998 25910 25050
rect 25962 24998 25974 25050
rect 26026 24998 28336 25050
rect 1104 24976 28336 24998
rect 1104 24506 28336 24528
rect 1104 24454 3282 24506
rect 3334 24454 3346 24506
rect 3398 24454 3410 24506
rect 3462 24454 3474 24506
rect 3526 24454 6282 24506
rect 6334 24454 6346 24506
rect 6398 24454 6410 24506
rect 6462 24454 6474 24506
rect 6526 24454 9282 24506
rect 9334 24454 9346 24506
rect 9398 24454 9410 24506
rect 9462 24454 9474 24506
rect 9526 24454 12282 24506
rect 12334 24454 12346 24506
rect 12398 24454 12410 24506
rect 12462 24454 12474 24506
rect 12526 24454 15282 24506
rect 15334 24454 15346 24506
rect 15398 24454 15410 24506
rect 15462 24454 15474 24506
rect 15526 24454 18282 24506
rect 18334 24454 18346 24506
rect 18398 24454 18410 24506
rect 18462 24454 18474 24506
rect 18526 24454 21282 24506
rect 21334 24454 21346 24506
rect 21398 24454 21410 24506
rect 21462 24454 21474 24506
rect 21526 24454 24282 24506
rect 24334 24454 24346 24506
rect 24398 24454 24410 24506
rect 24462 24454 24474 24506
rect 24526 24454 27282 24506
rect 27334 24454 27346 24506
rect 27398 24454 27410 24506
rect 27462 24454 27474 24506
rect 27526 24454 28336 24506
rect 1104 24432 28336 24454
rect 1104 23962 28336 23984
rect 1104 23910 1782 23962
rect 1834 23910 1846 23962
rect 1898 23910 1910 23962
rect 1962 23910 1974 23962
rect 2026 23910 4782 23962
rect 4834 23910 4846 23962
rect 4898 23910 4910 23962
rect 4962 23910 4974 23962
rect 5026 23910 7782 23962
rect 7834 23910 7846 23962
rect 7898 23910 7910 23962
rect 7962 23910 7974 23962
rect 8026 23910 10782 23962
rect 10834 23910 10846 23962
rect 10898 23910 10910 23962
rect 10962 23910 10974 23962
rect 11026 23910 13782 23962
rect 13834 23910 13846 23962
rect 13898 23910 13910 23962
rect 13962 23910 13974 23962
rect 14026 23910 16782 23962
rect 16834 23910 16846 23962
rect 16898 23910 16910 23962
rect 16962 23910 16974 23962
rect 17026 23910 19782 23962
rect 19834 23910 19846 23962
rect 19898 23910 19910 23962
rect 19962 23910 19974 23962
rect 20026 23910 22782 23962
rect 22834 23910 22846 23962
rect 22898 23910 22910 23962
rect 22962 23910 22974 23962
rect 23026 23910 25782 23962
rect 25834 23910 25846 23962
rect 25898 23910 25910 23962
rect 25962 23910 25974 23962
rect 26026 23910 28336 23962
rect 1104 23888 28336 23910
rect 1104 23418 28336 23440
rect 1104 23366 3282 23418
rect 3334 23366 3346 23418
rect 3398 23366 3410 23418
rect 3462 23366 3474 23418
rect 3526 23366 6282 23418
rect 6334 23366 6346 23418
rect 6398 23366 6410 23418
rect 6462 23366 6474 23418
rect 6526 23366 9282 23418
rect 9334 23366 9346 23418
rect 9398 23366 9410 23418
rect 9462 23366 9474 23418
rect 9526 23366 12282 23418
rect 12334 23366 12346 23418
rect 12398 23366 12410 23418
rect 12462 23366 12474 23418
rect 12526 23366 15282 23418
rect 15334 23366 15346 23418
rect 15398 23366 15410 23418
rect 15462 23366 15474 23418
rect 15526 23366 18282 23418
rect 18334 23366 18346 23418
rect 18398 23366 18410 23418
rect 18462 23366 18474 23418
rect 18526 23366 21282 23418
rect 21334 23366 21346 23418
rect 21398 23366 21410 23418
rect 21462 23366 21474 23418
rect 21526 23366 24282 23418
rect 24334 23366 24346 23418
rect 24398 23366 24410 23418
rect 24462 23366 24474 23418
rect 24526 23366 27282 23418
rect 27334 23366 27346 23418
rect 27398 23366 27410 23418
rect 27462 23366 27474 23418
rect 27526 23366 28336 23418
rect 1104 23344 28336 23366
rect 1104 22874 28336 22896
rect 1104 22822 1782 22874
rect 1834 22822 1846 22874
rect 1898 22822 1910 22874
rect 1962 22822 1974 22874
rect 2026 22822 4782 22874
rect 4834 22822 4846 22874
rect 4898 22822 4910 22874
rect 4962 22822 4974 22874
rect 5026 22822 7782 22874
rect 7834 22822 7846 22874
rect 7898 22822 7910 22874
rect 7962 22822 7974 22874
rect 8026 22822 10782 22874
rect 10834 22822 10846 22874
rect 10898 22822 10910 22874
rect 10962 22822 10974 22874
rect 11026 22822 13782 22874
rect 13834 22822 13846 22874
rect 13898 22822 13910 22874
rect 13962 22822 13974 22874
rect 14026 22822 16782 22874
rect 16834 22822 16846 22874
rect 16898 22822 16910 22874
rect 16962 22822 16974 22874
rect 17026 22822 19782 22874
rect 19834 22822 19846 22874
rect 19898 22822 19910 22874
rect 19962 22822 19974 22874
rect 20026 22822 22782 22874
rect 22834 22822 22846 22874
rect 22898 22822 22910 22874
rect 22962 22822 22974 22874
rect 23026 22822 25782 22874
rect 25834 22822 25846 22874
rect 25898 22822 25910 22874
rect 25962 22822 25974 22874
rect 26026 22822 28336 22874
rect 1104 22800 28336 22822
rect 1104 22330 28336 22352
rect 1104 22278 3282 22330
rect 3334 22278 3346 22330
rect 3398 22278 3410 22330
rect 3462 22278 3474 22330
rect 3526 22278 6282 22330
rect 6334 22278 6346 22330
rect 6398 22278 6410 22330
rect 6462 22278 6474 22330
rect 6526 22278 9282 22330
rect 9334 22278 9346 22330
rect 9398 22278 9410 22330
rect 9462 22278 9474 22330
rect 9526 22278 12282 22330
rect 12334 22278 12346 22330
rect 12398 22278 12410 22330
rect 12462 22278 12474 22330
rect 12526 22278 15282 22330
rect 15334 22278 15346 22330
rect 15398 22278 15410 22330
rect 15462 22278 15474 22330
rect 15526 22278 18282 22330
rect 18334 22278 18346 22330
rect 18398 22278 18410 22330
rect 18462 22278 18474 22330
rect 18526 22278 21282 22330
rect 21334 22278 21346 22330
rect 21398 22278 21410 22330
rect 21462 22278 21474 22330
rect 21526 22278 24282 22330
rect 24334 22278 24346 22330
rect 24398 22278 24410 22330
rect 24462 22278 24474 22330
rect 24526 22278 27282 22330
rect 27334 22278 27346 22330
rect 27398 22278 27410 22330
rect 27462 22278 27474 22330
rect 27526 22278 28336 22330
rect 1104 22256 28336 22278
rect 1104 21786 28336 21808
rect 1104 21734 1782 21786
rect 1834 21734 1846 21786
rect 1898 21734 1910 21786
rect 1962 21734 1974 21786
rect 2026 21734 4782 21786
rect 4834 21734 4846 21786
rect 4898 21734 4910 21786
rect 4962 21734 4974 21786
rect 5026 21734 7782 21786
rect 7834 21734 7846 21786
rect 7898 21734 7910 21786
rect 7962 21734 7974 21786
rect 8026 21734 10782 21786
rect 10834 21734 10846 21786
rect 10898 21734 10910 21786
rect 10962 21734 10974 21786
rect 11026 21734 13782 21786
rect 13834 21734 13846 21786
rect 13898 21734 13910 21786
rect 13962 21734 13974 21786
rect 14026 21734 16782 21786
rect 16834 21734 16846 21786
rect 16898 21734 16910 21786
rect 16962 21734 16974 21786
rect 17026 21734 19782 21786
rect 19834 21734 19846 21786
rect 19898 21734 19910 21786
rect 19962 21734 19974 21786
rect 20026 21734 22782 21786
rect 22834 21734 22846 21786
rect 22898 21734 22910 21786
rect 22962 21734 22974 21786
rect 23026 21734 25782 21786
rect 25834 21734 25846 21786
rect 25898 21734 25910 21786
rect 25962 21734 25974 21786
rect 26026 21734 28336 21786
rect 1104 21712 28336 21734
rect 1104 21242 28336 21264
rect 1104 21190 3282 21242
rect 3334 21190 3346 21242
rect 3398 21190 3410 21242
rect 3462 21190 3474 21242
rect 3526 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 6410 21242
rect 6462 21190 6474 21242
rect 6526 21190 9282 21242
rect 9334 21190 9346 21242
rect 9398 21190 9410 21242
rect 9462 21190 9474 21242
rect 9526 21190 12282 21242
rect 12334 21190 12346 21242
rect 12398 21190 12410 21242
rect 12462 21190 12474 21242
rect 12526 21190 15282 21242
rect 15334 21190 15346 21242
rect 15398 21190 15410 21242
rect 15462 21190 15474 21242
rect 15526 21190 18282 21242
rect 18334 21190 18346 21242
rect 18398 21190 18410 21242
rect 18462 21190 18474 21242
rect 18526 21190 21282 21242
rect 21334 21190 21346 21242
rect 21398 21190 21410 21242
rect 21462 21190 21474 21242
rect 21526 21190 24282 21242
rect 24334 21190 24346 21242
rect 24398 21190 24410 21242
rect 24462 21190 24474 21242
rect 24526 21190 27282 21242
rect 27334 21190 27346 21242
rect 27398 21190 27410 21242
rect 27462 21190 27474 21242
rect 27526 21190 28336 21242
rect 1104 21168 28336 21190
rect 1104 20698 28336 20720
rect 1104 20646 1782 20698
rect 1834 20646 1846 20698
rect 1898 20646 1910 20698
rect 1962 20646 1974 20698
rect 2026 20646 4782 20698
rect 4834 20646 4846 20698
rect 4898 20646 4910 20698
rect 4962 20646 4974 20698
rect 5026 20646 7782 20698
rect 7834 20646 7846 20698
rect 7898 20646 7910 20698
rect 7962 20646 7974 20698
rect 8026 20646 10782 20698
rect 10834 20646 10846 20698
rect 10898 20646 10910 20698
rect 10962 20646 10974 20698
rect 11026 20646 13782 20698
rect 13834 20646 13846 20698
rect 13898 20646 13910 20698
rect 13962 20646 13974 20698
rect 14026 20646 16782 20698
rect 16834 20646 16846 20698
rect 16898 20646 16910 20698
rect 16962 20646 16974 20698
rect 17026 20646 19782 20698
rect 19834 20646 19846 20698
rect 19898 20646 19910 20698
rect 19962 20646 19974 20698
rect 20026 20646 22782 20698
rect 22834 20646 22846 20698
rect 22898 20646 22910 20698
rect 22962 20646 22974 20698
rect 23026 20646 25782 20698
rect 25834 20646 25846 20698
rect 25898 20646 25910 20698
rect 25962 20646 25974 20698
rect 26026 20646 28336 20698
rect 1104 20624 28336 20646
rect 1104 20154 28336 20176
rect 1104 20102 3282 20154
rect 3334 20102 3346 20154
rect 3398 20102 3410 20154
rect 3462 20102 3474 20154
rect 3526 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 6410 20154
rect 6462 20102 6474 20154
rect 6526 20102 9282 20154
rect 9334 20102 9346 20154
rect 9398 20102 9410 20154
rect 9462 20102 9474 20154
rect 9526 20102 12282 20154
rect 12334 20102 12346 20154
rect 12398 20102 12410 20154
rect 12462 20102 12474 20154
rect 12526 20102 15282 20154
rect 15334 20102 15346 20154
rect 15398 20102 15410 20154
rect 15462 20102 15474 20154
rect 15526 20102 18282 20154
rect 18334 20102 18346 20154
rect 18398 20102 18410 20154
rect 18462 20102 18474 20154
rect 18526 20102 21282 20154
rect 21334 20102 21346 20154
rect 21398 20102 21410 20154
rect 21462 20102 21474 20154
rect 21526 20102 24282 20154
rect 24334 20102 24346 20154
rect 24398 20102 24410 20154
rect 24462 20102 24474 20154
rect 24526 20102 27282 20154
rect 27334 20102 27346 20154
rect 27398 20102 27410 20154
rect 27462 20102 27474 20154
rect 27526 20102 28336 20154
rect 1104 20080 28336 20102
rect 1104 19610 28336 19632
rect 1104 19558 1782 19610
rect 1834 19558 1846 19610
rect 1898 19558 1910 19610
rect 1962 19558 1974 19610
rect 2026 19558 4782 19610
rect 4834 19558 4846 19610
rect 4898 19558 4910 19610
rect 4962 19558 4974 19610
rect 5026 19558 7782 19610
rect 7834 19558 7846 19610
rect 7898 19558 7910 19610
rect 7962 19558 7974 19610
rect 8026 19558 10782 19610
rect 10834 19558 10846 19610
rect 10898 19558 10910 19610
rect 10962 19558 10974 19610
rect 11026 19558 13782 19610
rect 13834 19558 13846 19610
rect 13898 19558 13910 19610
rect 13962 19558 13974 19610
rect 14026 19558 16782 19610
rect 16834 19558 16846 19610
rect 16898 19558 16910 19610
rect 16962 19558 16974 19610
rect 17026 19558 19782 19610
rect 19834 19558 19846 19610
rect 19898 19558 19910 19610
rect 19962 19558 19974 19610
rect 20026 19558 22782 19610
rect 22834 19558 22846 19610
rect 22898 19558 22910 19610
rect 22962 19558 22974 19610
rect 23026 19558 25782 19610
rect 25834 19558 25846 19610
rect 25898 19558 25910 19610
rect 25962 19558 25974 19610
rect 26026 19558 28336 19610
rect 1104 19536 28336 19558
rect 1104 19066 28336 19088
rect 1104 19014 3282 19066
rect 3334 19014 3346 19066
rect 3398 19014 3410 19066
rect 3462 19014 3474 19066
rect 3526 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 6410 19066
rect 6462 19014 6474 19066
rect 6526 19014 9282 19066
rect 9334 19014 9346 19066
rect 9398 19014 9410 19066
rect 9462 19014 9474 19066
rect 9526 19014 12282 19066
rect 12334 19014 12346 19066
rect 12398 19014 12410 19066
rect 12462 19014 12474 19066
rect 12526 19014 15282 19066
rect 15334 19014 15346 19066
rect 15398 19014 15410 19066
rect 15462 19014 15474 19066
rect 15526 19014 18282 19066
rect 18334 19014 18346 19066
rect 18398 19014 18410 19066
rect 18462 19014 18474 19066
rect 18526 19014 21282 19066
rect 21334 19014 21346 19066
rect 21398 19014 21410 19066
rect 21462 19014 21474 19066
rect 21526 19014 24282 19066
rect 24334 19014 24346 19066
rect 24398 19014 24410 19066
rect 24462 19014 24474 19066
rect 24526 19014 27282 19066
rect 27334 19014 27346 19066
rect 27398 19014 27410 19066
rect 27462 19014 27474 19066
rect 27526 19014 28336 19066
rect 1104 18992 28336 19014
rect 1104 18522 28336 18544
rect 1104 18470 1782 18522
rect 1834 18470 1846 18522
rect 1898 18470 1910 18522
rect 1962 18470 1974 18522
rect 2026 18470 4782 18522
rect 4834 18470 4846 18522
rect 4898 18470 4910 18522
rect 4962 18470 4974 18522
rect 5026 18470 7782 18522
rect 7834 18470 7846 18522
rect 7898 18470 7910 18522
rect 7962 18470 7974 18522
rect 8026 18470 10782 18522
rect 10834 18470 10846 18522
rect 10898 18470 10910 18522
rect 10962 18470 10974 18522
rect 11026 18470 13782 18522
rect 13834 18470 13846 18522
rect 13898 18470 13910 18522
rect 13962 18470 13974 18522
rect 14026 18470 16782 18522
rect 16834 18470 16846 18522
rect 16898 18470 16910 18522
rect 16962 18470 16974 18522
rect 17026 18470 19782 18522
rect 19834 18470 19846 18522
rect 19898 18470 19910 18522
rect 19962 18470 19974 18522
rect 20026 18470 22782 18522
rect 22834 18470 22846 18522
rect 22898 18470 22910 18522
rect 22962 18470 22974 18522
rect 23026 18470 25782 18522
rect 25834 18470 25846 18522
rect 25898 18470 25910 18522
rect 25962 18470 25974 18522
rect 26026 18470 28336 18522
rect 1104 18448 28336 18470
rect 1104 17978 28336 18000
rect 1104 17926 3282 17978
rect 3334 17926 3346 17978
rect 3398 17926 3410 17978
rect 3462 17926 3474 17978
rect 3526 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 6410 17978
rect 6462 17926 6474 17978
rect 6526 17926 9282 17978
rect 9334 17926 9346 17978
rect 9398 17926 9410 17978
rect 9462 17926 9474 17978
rect 9526 17926 12282 17978
rect 12334 17926 12346 17978
rect 12398 17926 12410 17978
rect 12462 17926 12474 17978
rect 12526 17926 15282 17978
rect 15334 17926 15346 17978
rect 15398 17926 15410 17978
rect 15462 17926 15474 17978
rect 15526 17926 18282 17978
rect 18334 17926 18346 17978
rect 18398 17926 18410 17978
rect 18462 17926 18474 17978
rect 18526 17926 21282 17978
rect 21334 17926 21346 17978
rect 21398 17926 21410 17978
rect 21462 17926 21474 17978
rect 21526 17926 24282 17978
rect 24334 17926 24346 17978
rect 24398 17926 24410 17978
rect 24462 17926 24474 17978
rect 24526 17926 27282 17978
rect 27334 17926 27346 17978
rect 27398 17926 27410 17978
rect 27462 17926 27474 17978
rect 27526 17926 28336 17978
rect 1104 17904 28336 17926
rect 1104 17434 28336 17456
rect 1104 17382 1782 17434
rect 1834 17382 1846 17434
rect 1898 17382 1910 17434
rect 1962 17382 1974 17434
rect 2026 17382 4782 17434
rect 4834 17382 4846 17434
rect 4898 17382 4910 17434
rect 4962 17382 4974 17434
rect 5026 17382 7782 17434
rect 7834 17382 7846 17434
rect 7898 17382 7910 17434
rect 7962 17382 7974 17434
rect 8026 17382 10782 17434
rect 10834 17382 10846 17434
rect 10898 17382 10910 17434
rect 10962 17382 10974 17434
rect 11026 17382 13782 17434
rect 13834 17382 13846 17434
rect 13898 17382 13910 17434
rect 13962 17382 13974 17434
rect 14026 17382 16782 17434
rect 16834 17382 16846 17434
rect 16898 17382 16910 17434
rect 16962 17382 16974 17434
rect 17026 17382 19782 17434
rect 19834 17382 19846 17434
rect 19898 17382 19910 17434
rect 19962 17382 19974 17434
rect 20026 17382 22782 17434
rect 22834 17382 22846 17434
rect 22898 17382 22910 17434
rect 22962 17382 22974 17434
rect 23026 17382 25782 17434
rect 25834 17382 25846 17434
rect 25898 17382 25910 17434
rect 25962 17382 25974 17434
rect 26026 17382 28336 17434
rect 1104 17360 28336 17382
rect 1104 16890 28336 16912
rect 1104 16838 3282 16890
rect 3334 16838 3346 16890
rect 3398 16838 3410 16890
rect 3462 16838 3474 16890
rect 3526 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 6410 16890
rect 6462 16838 6474 16890
rect 6526 16838 9282 16890
rect 9334 16838 9346 16890
rect 9398 16838 9410 16890
rect 9462 16838 9474 16890
rect 9526 16838 12282 16890
rect 12334 16838 12346 16890
rect 12398 16838 12410 16890
rect 12462 16838 12474 16890
rect 12526 16838 15282 16890
rect 15334 16838 15346 16890
rect 15398 16838 15410 16890
rect 15462 16838 15474 16890
rect 15526 16838 18282 16890
rect 18334 16838 18346 16890
rect 18398 16838 18410 16890
rect 18462 16838 18474 16890
rect 18526 16838 21282 16890
rect 21334 16838 21346 16890
rect 21398 16838 21410 16890
rect 21462 16838 21474 16890
rect 21526 16838 24282 16890
rect 24334 16838 24346 16890
rect 24398 16838 24410 16890
rect 24462 16838 24474 16890
rect 24526 16838 27282 16890
rect 27334 16838 27346 16890
rect 27398 16838 27410 16890
rect 27462 16838 27474 16890
rect 27526 16838 28336 16890
rect 1104 16816 28336 16838
rect 14090 16572 14096 16584
rect 14051 16544 14096 16572
rect 14090 16532 14096 16544
rect 14148 16532 14154 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15620 16544 15669 16572
rect 15620 16532 15626 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 15473 16507 15531 16513
rect 15473 16473 15485 16507
rect 15519 16504 15531 16507
rect 15746 16504 15752 16516
rect 15519 16476 15752 16504
rect 15519 16473 15531 16476
rect 15473 16467 15531 16473
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 16025 16507 16083 16513
rect 16025 16473 16037 16507
rect 16071 16504 16083 16507
rect 16482 16504 16488 16516
rect 16071 16476 16488 16504
rect 16071 16473 16083 16476
rect 16025 16467 16083 16473
rect 16482 16464 16488 16476
rect 16540 16464 16546 16516
rect 14274 16436 14280 16448
rect 14235 16408 14280 16436
rect 14274 16396 14280 16408
rect 14332 16436 14338 16448
rect 14918 16436 14924 16448
rect 14332 16408 14924 16436
rect 14332 16396 14338 16408
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 1104 16346 28336 16368
rect 1104 16294 1782 16346
rect 1834 16294 1846 16346
rect 1898 16294 1910 16346
rect 1962 16294 1974 16346
rect 2026 16294 4782 16346
rect 4834 16294 4846 16346
rect 4898 16294 4910 16346
rect 4962 16294 4974 16346
rect 5026 16294 7782 16346
rect 7834 16294 7846 16346
rect 7898 16294 7910 16346
rect 7962 16294 7974 16346
rect 8026 16294 10782 16346
rect 10834 16294 10846 16346
rect 10898 16294 10910 16346
rect 10962 16294 10974 16346
rect 11026 16294 13782 16346
rect 13834 16294 13846 16346
rect 13898 16294 13910 16346
rect 13962 16294 13974 16346
rect 14026 16294 16782 16346
rect 16834 16294 16846 16346
rect 16898 16294 16910 16346
rect 16962 16294 16974 16346
rect 17026 16294 19782 16346
rect 19834 16294 19846 16346
rect 19898 16294 19910 16346
rect 19962 16294 19974 16346
rect 20026 16294 22782 16346
rect 22834 16294 22846 16346
rect 22898 16294 22910 16346
rect 22962 16294 22974 16346
rect 23026 16294 25782 16346
rect 25834 16294 25846 16346
rect 25898 16294 25910 16346
rect 25962 16294 25974 16346
rect 26026 16294 28336 16346
rect 1104 16272 28336 16294
rect 14918 16124 14924 16176
rect 14976 16124 14982 16176
rect 14182 16028 14188 16040
rect 14143 16000 14188 16028
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 14550 16028 14556 16040
rect 14507 16000 14556 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15712 16000 16221 16028
rect 15712 15988 15718 16000
rect 16209 15997 16221 16000
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 15562 15920 15568 15972
rect 15620 15960 15626 15972
rect 16485 15963 16543 15969
rect 16485 15960 16497 15963
rect 15620 15932 16497 15960
rect 15620 15920 15626 15932
rect 16485 15929 16497 15932
rect 16531 15929 16543 15963
rect 16485 15923 16543 15929
rect 13909 15895 13967 15901
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 14090 15892 14096 15904
rect 13955 15864 14096 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 16574 15852 16580 15904
rect 16632 15892 16638 15904
rect 16853 15895 16911 15901
rect 16853 15892 16865 15895
rect 16632 15864 16865 15892
rect 16632 15852 16638 15864
rect 16853 15861 16865 15864
rect 16899 15861 16911 15895
rect 17310 15892 17316 15904
rect 17271 15864 17316 15892
rect 16853 15855 16911 15861
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 1104 15802 28336 15824
rect 1104 15750 3282 15802
rect 3334 15750 3346 15802
rect 3398 15750 3410 15802
rect 3462 15750 3474 15802
rect 3526 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 6410 15802
rect 6462 15750 6474 15802
rect 6526 15750 9282 15802
rect 9334 15750 9346 15802
rect 9398 15750 9410 15802
rect 9462 15750 9474 15802
rect 9526 15750 12282 15802
rect 12334 15750 12346 15802
rect 12398 15750 12410 15802
rect 12462 15750 12474 15802
rect 12526 15750 15282 15802
rect 15334 15750 15346 15802
rect 15398 15750 15410 15802
rect 15462 15750 15474 15802
rect 15526 15750 18282 15802
rect 18334 15750 18346 15802
rect 18398 15750 18410 15802
rect 18462 15750 18474 15802
rect 18526 15750 21282 15802
rect 21334 15750 21346 15802
rect 21398 15750 21410 15802
rect 21462 15750 21474 15802
rect 21526 15750 24282 15802
rect 24334 15750 24346 15802
rect 24398 15750 24410 15802
rect 24462 15750 24474 15802
rect 24526 15750 27282 15802
rect 27334 15750 27346 15802
rect 27398 15750 27410 15802
rect 27462 15750 27474 15802
rect 27526 15750 28336 15802
rect 1104 15728 28336 15750
rect 13909 15691 13967 15697
rect 13909 15657 13921 15691
rect 13955 15688 13967 15691
rect 14274 15688 14280 15700
rect 13955 15660 14280 15688
rect 13955 15657 13967 15660
rect 13909 15651 13967 15657
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 15746 15620 15752 15632
rect 15659 15592 15752 15620
rect 12710 15484 12716 15496
rect 12671 15456 12716 15484
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15672 15493 15700 15592
rect 15746 15580 15752 15592
rect 15804 15620 15810 15632
rect 16574 15620 16580 15632
rect 15804 15592 16580 15620
rect 15804 15580 15810 15592
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 16761 15555 16819 15561
rect 16761 15552 16773 15555
rect 16264 15524 16773 15552
rect 16264 15512 16270 15524
rect 16761 15521 16773 15524
rect 16807 15521 16819 15555
rect 16761 15515 16819 15521
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15436 15456 15669 15484
rect 15436 15444 15442 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 15657 15447 15715 15453
rect 16408 15456 17233 15484
rect 15470 15416 15476 15428
rect 15431 15388 15476 15416
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 16022 15416 16028 15428
rect 15983 15388 16028 15416
rect 16022 15376 16028 15388
rect 16080 15376 16086 15428
rect 16408 15360 16436 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17310 15444 17316 15496
rect 17368 15484 17374 15496
rect 17405 15487 17463 15493
rect 17405 15484 17417 15487
rect 17368 15456 17417 15484
rect 17368 15444 17374 15456
rect 17405 15453 17417 15456
rect 17451 15453 17463 15487
rect 17770 15484 17776 15496
rect 17731 15456 17776 15484
rect 17405 15447 17463 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18138 15484 18144 15496
rect 18003 15456 18144 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 18564 15456 19441 15484
rect 18564 15444 18570 15456
rect 19429 15453 19441 15456
rect 19475 15484 19487 15487
rect 20530 15484 20536 15496
rect 19475 15456 20536 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 12894 15348 12900 15360
rect 12855 15320 12900 15348
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13262 15348 13268 15360
rect 13223 15320 13268 15348
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 14182 15348 14188 15360
rect 14143 15320 14188 15348
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14642 15348 14648 15360
rect 14603 15320 14648 15348
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 16390 15348 16396 15360
rect 16351 15320 16396 15348
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 18509 15351 18567 15357
rect 18509 15317 18521 15351
rect 18555 15348 18567 15351
rect 18782 15348 18788 15360
rect 18555 15320 18788 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 19061 15351 19119 15357
rect 19061 15317 19073 15351
rect 19107 15348 19119 15351
rect 19150 15348 19156 15360
rect 19107 15320 19156 15348
rect 19107 15317 19119 15320
rect 19061 15311 19119 15317
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 1104 15258 28336 15280
rect 1104 15206 1782 15258
rect 1834 15206 1846 15258
rect 1898 15206 1910 15258
rect 1962 15206 1974 15258
rect 2026 15206 4782 15258
rect 4834 15206 4846 15258
rect 4898 15206 4910 15258
rect 4962 15206 4974 15258
rect 5026 15206 7782 15258
rect 7834 15206 7846 15258
rect 7898 15206 7910 15258
rect 7962 15206 7974 15258
rect 8026 15206 10782 15258
rect 10834 15206 10846 15258
rect 10898 15206 10910 15258
rect 10962 15206 10974 15258
rect 11026 15206 13782 15258
rect 13834 15206 13846 15258
rect 13898 15206 13910 15258
rect 13962 15206 13974 15258
rect 14026 15206 16782 15258
rect 16834 15206 16846 15258
rect 16898 15206 16910 15258
rect 16962 15206 16974 15258
rect 17026 15206 19782 15258
rect 19834 15206 19846 15258
rect 19898 15206 19910 15258
rect 19962 15206 19974 15258
rect 20026 15206 22782 15258
rect 22834 15206 22846 15258
rect 22898 15206 22910 15258
rect 22962 15206 22974 15258
rect 23026 15206 25782 15258
rect 25834 15206 25846 15258
rect 25898 15206 25910 15258
rect 25962 15206 25974 15258
rect 26026 15206 28336 15258
rect 1104 15184 28336 15206
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12768 15116 12817 15144
rect 12768 15104 12774 15116
rect 12805 15113 12817 15116
rect 12851 15144 12863 15147
rect 14090 15144 14096 15156
rect 12851 15116 14096 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 14090 15104 14096 15116
rect 14148 15144 14154 15156
rect 15378 15144 15384 15156
rect 14148 15116 14228 15144
rect 15339 15116 15384 15144
rect 14148 15104 14154 15116
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 13814 15008 13820 15020
rect 13320 14980 13820 15008
rect 13320 14968 13326 14980
rect 13814 14968 13820 14980
rect 13872 15008 13878 15020
rect 13872 14980 13917 15008
rect 13872 14968 13878 14980
rect 14200 14872 14228 15116
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 16301 15147 16359 15153
rect 16301 15113 16313 15147
rect 16347 15144 16359 15147
rect 17770 15144 17776 15156
rect 16347 15116 17776 15144
rect 16347 15113 16359 15116
rect 16301 15107 16359 15113
rect 17770 15104 17776 15116
rect 17828 15144 17834 15156
rect 18874 15144 18880 15156
rect 17828 15116 18880 15144
rect 17828 15104 17834 15116
rect 14645 15079 14703 15085
rect 14645 15045 14657 15079
rect 14691 15076 14703 15079
rect 14826 15076 14832 15088
rect 14691 15048 14832 15076
rect 14691 15045 14703 15048
rect 14645 15039 14703 15045
rect 14826 15036 14832 15048
rect 14884 15076 14890 15088
rect 15470 15076 15476 15088
rect 14884 15048 15476 15076
rect 14884 15036 14890 15048
rect 15470 15036 15476 15048
rect 15528 15076 15534 15088
rect 17129 15079 17187 15085
rect 15528 15048 16712 15076
rect 15528 15036 15534 15048
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14550 15008 14556 15020
rect 14323 14980 14556 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 14550 14968 14556 14980
rect 14608 15008 14614 15020
rect 15010 15008 15016 15020
rect 14608 14980 15016 15008
rect 14608 14968 14614 14980
rect 15010 14968 15016 14980
rect 15068 15008 15074 15020
rect 15565 15011 15623 15017
rect 15565 15008 15577 15011
rect 15068 14980 15577 15008
rect 15068 14968 15074 14980
rect 15565 14977 15577 14980
rect 15611 15008 15623 15011
rect 15654 15008 15660 15020
rect 15611 14980 15660 15008
rect 15611 14977 15623 14980
rect 15565 14971 15623 14977
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 16574 15008 16580 15020
rect 16535 14980 16580 15008
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16684 15017 16712 15048
rect 17129 15045 17141 15079
rect 17175 15076 17187 15079
rect 17310 15076 17316 15088
rect 17175 15048 17316 15076
rect 17175 15045 17187 15048
rect 17129 15039 17187 15045
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 17494 15036 17500 15088
rect 17552 15076 17558 15088
rect 18506 15076 18512 15088
rect 17552 15048 18512 15076
rect 17552 15036 17558 15048
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 18800 15085 18828 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 18785 15079 18843 15085
rect 18785 15045 18797 15079
rect 18831 15045 18843 15079
rect 18785 15039 18843 15045
rect 21174 15036 21180 15088
rect 21232 15036 21238 15088
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 17512 15008 17540 15036
rect 16715 14980 17540 15008
rect 19429 15011 19487 15017
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 19429 14977 19441 15011
rect 19475 15008 19487 15011
rect 19475 14980 19932 15008
rect 19475 14977 19487 14980
rect 19429 14971 19487 14977
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19444 14940 19472 14971
rect 18840 14912 19472 14940
rect 18840 14900 18846 14912
rect 19426 14872 19432 14884
rect 14200 14844 19432 14872
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 13630 14804 13636 14816
rect 13591 14776 13636 14804
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 17497 14807 17555 14813
rect 17497 14773 17509 14807
rect 17543 14804 17555 14807
rect 18138 14804 18144 14816
rect 17543 14776 18144 14804
rect 17543 14773 17555 14776
rect 17497 14767 17555 14773
rect 18138 14764 18144 14776
rect 18196 14764 18202 14816
rect 19904 14813 19932 14980
rect 20346 14940 20352 14952
rect 20307 14912 20352 14940
rect 20346 14900 20352 14912
rect 20404 14900 20410 14952
rect 20622 14940 20628 14952
rect 20583 14912 20628 14940
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 22373 14943 22431 14949
rect 22373 14909 22385 14943
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 19889 14807 19947 14813
rect 19889 14773 19901 14807
rect 19935 14804 19947 14807
rect 20714 14804 20720 14816
rect 19935 14776 20720 14804
rect 19935 14773 19947 14776
rect 19889 14767 19947 14773
rect 20714 14764 20720 14776
rect 20772 14804 20778 14816
rect 22388 14804 22416 14903
rect 20772 14776 22416 14804
rect 20772 14764 20778 14776
rect 1104 14714 28336 14736
rect 1104 14662 3282 14714
rect 3334 14662 3346 14714
rect 3398 14662 3410 14714
rect 3462 14662 3474 14714
rect 3526 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 6410 14714
rect 6462 14662 6474 14714
rect 6526 14662 9282 14714
rect 9334 14662 9346 14714
rect 9398 14662 9410 14714
rect 9462 14662 9474 14714
rect 9526 14662 12282 14714
rect 12334 14662 12346 14714
rect 12398 14662 12410 14714
rect 12462 14662 12474 14714
rect 12526 14662 15282 14714
rect 15334 14662 15346 14714
rect 15398 14662 15410 14714
rect 15462 14662 15474 14714
rect 15526 14662 18282 14714
rect 18334 14662 18346 14714
rect 18398 14662 18410 14714
rect 18462 14662 18474 14714
rect 18526 14662 21282 14714
rect 21334 14662 21346 14714
rect 21398 14662 21410 14714
rect 21462 14662 21474 14714
rect 21526 14662 24282 14714
rect 24334 14662 24346 14714
rect 24398 14662 24410 14714
rect 24462 14662 24474 14714
rect 24526 14662 27282 14714
rect 27334 14662 27346 14714
rect 27398 14662 27410 14714
rect 27462 14662 27474 14714
rect 27526 14662 28336 14714
rect 1104 14640 28336 14662
rect 14550 14600 14556 14612
rect 14511 14572 14556 14600
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 14921 14603 14979 14609
rect 14921 14569 14933 14603
rect 14967 14600 14979 14603
rect 15102 14600 15108 14612
rect 14967 14572 15108 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 15102 14560 15108 14572
rect 15160 14600 15166 14612
rect 16574 14600 16580 14612
rect 15160 14572 16580 14600
rect 15160 14560 15166 14572
rect 16574 14560 16580 14572
rect 16632 14600 16638 14612
rect 17405 14603 17463 14609
rect 17405 14600 17417 14603
rect 16632 14572 17417 14600
rect 16632 14560 16638 14572
rect 17405 14569 17417 14572
rect 17451 14569 17463 14603
rect 17405 14563 17463 14569
rect 21174 14560 21180 14612
rect 21232 14600 21238 14612
rect 21361 14603 21419 14609
rect 21361 14600 21373 14603
rect 21232 14572 21373 14600
rect 21232 14560 21238 14572
rect 21361 14569 21373 14572
rect 21407 14600 21419 14603
rect 21637 14603 21695 14609
rect 21637 14600 21649 14603
rect 21407 14572 21649 14600
rect 21407 14569 21419 14572
rect 21361 14563 21419 14569
rect 21637 14569 21649 14572
rect 21683 14569 21695 14603
rect 21637 14563 21695 14569
rect 14642 14492 14648 14544
rect 14700 14532 14706 14544
rect 16485 14535 16543 14541
rect 16485 14532 16497 14535
rect 14700 14504 16497 14532
rect 14700 14492 14706 14504
rect 16485 14501 16497 14504
rect 16531 14501 16543 14535
rect 16485 14495 16543 14501
rect 17129 14535 17187 14541
rect 17129 14501 17141 14535
rect 17175 14532 17187 14535
rect 17494 14532 17500 14544
rect 17175 14504 17500 14532
rect 17175 14501 17187 14504
rect 17129 14495 17187 14501
rect 17494 14492 17500 14504
rect 17552 14492 17558 14544
rect 11882 14464 11888 14476
rect 11795 14436 11888 14464
rect 11882 14424 11888 14436
rect 11940 14464 11946 14476
rect 14182 14464 14188 14476
rect 11940 14436 14188 14464
rect 11940 14424 11946 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 18616 14436 18920 14464
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 15930 14396 15936 14408
rect 15887 14368 15936 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16206 14396 16212 14408
rect 16167 14368 16212 14396
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 16482 14396 16488 14408
rect 16443 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 18616 14405 18644 14436
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 17184 14368 18245 14396
rect 17184 14356 17190 14368
rect 18233 14365 18245 14368
rect 18279 14396 18291 14399
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18279 14368 18613 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18782 14396 18788 14408
rect 18743 14368 18788 14396
rect 18601 14359 18659 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 18892 14396 18920 14436
rect 19242 14396 19248 14408
rect 18892 14368 19248 14396
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 12158 14328 12164 14340
rect 12119 14300 12164 14328
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 12894 14288 12900 14340
rect 12952 14288 12958 14340
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 13909 14331 13967 14337
rect 13909 14328 13921 14331
rect 13872 14300 13921 14328
rect 13872 14288 13878 14300
rect 13909 14297 13921 14300
rect 13955 14328 13967 14331
rect 14274 14328 14280 14340
rect 13955 14300 14280 14328
rect 13955 14297 13967 14300
rect 13909 14291 13967 14297
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 19352 14328 19380 14359
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 21174 14396 21180 14408
rect 19484 14368 21180 14396
rect 19484 14356 19490 14368
rect 21174 14356 21180 14368
rect 21232 14356 21238 14408
rect 17972 14300 19380 14328
rect 19889 14331 19947 14337
rect 17972 14272 18000 14300
rect 19889 14297 19901 14331
rect 19935 14328 19947 14331
rect 20622 14328 20628 14340
rect 19935 14300 20628 14328
rect 19935 14297 19947 14300
rect 19889 14291 19947 14297
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 17954 14260 17960 14272
rect 17915 14232 17960 14260
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 20346 14260 20352 14272
rect 20307 14232 20352 14260
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 1104 14170 28336 14192
rect 1104 14118 1782 14170
rect 1834 14118 1846 14170
rect 1898 14118 1910 14170
rect 1962 14118 1974 14170
rect 2026 14118 4782 14170
rect 4834 14118 4846 14170
rect 4898 14118 4910 14170
rect 4962 14118 4974 14170
rect 5026 14118 7782 14170
rect 7834 14118 7846 14170
rect 7898 14118 7910 14170
rect 7962 14118 7974 14170
rect 8026 14118 10782 14170
rect 10834 14118 10846 14170
rect 10898 14118 10910 14170
rect 10962 14118 10974 14170
rect 11026 14118 13782 14170
rect 13834 14118 13846 14170
rect 13898 14118 13910 14170
rect 13962 14118 13974 14170
rect 14026 14118 16782 14170
rect 16834 14118 16846 14170
rect 16898 14118 16910 14170
rect 16962 14118 16974 14170
rect 17026 14118 19782 14170
rect 19834 14118 19846 14170
rect 19898 14118 19910 14170
rect 19962 14118 19974 14170
rect 20026 14118 22782 14170
rect 22834 14118 22846 14170
rect 22898 14118 22910 14170
rect 22962 14118 22974 14170
rect 23026 14118 25782 14170
rect 25834 14118 25846 14170
rect 25898 14118 25910 14170
rect 25962 14118 25974 14170
rect 26026 14118 28336 14170
rect 1104 14096 28336 14118
rect 11609 14059 11667 14065
rect 11609 14025 11621 14059
rect 11655 14056 11667 14059
rect 12158 14056 12164 14068
rect 11655 14028 12164 14056
rect 11655 14025 11667 14028
rect 11609 14019 11667 14025
rect 12158 14016 12164 14028
rect 12216 14056 12222 14068
rect 14553 14059 14611 14065
rect 12216 14028 12664 14056
rect 12216 14016 12222 14028
rect 11882 13988 11888 14000
rect 11843 13960 11888 13988
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 12636 13997 12664 14028
rect 14553 14025 14565 14059
rect 14599 14056 14611 14059
rect 16206 14056 16212 14068
rect 14599 14028 16212 14056
rect 14599 14025 14611 14028
rect 14553 14019 14611 14025
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17052 14028 17693 14056
rect 17052 14000 17080 14028
rect 17681 14025 17693 14028
rect 17727 14056 17739 14059
rect 19150 14056 19156 14068
rect 17727 14028 19156 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19300 14028 19901 14056
rect 19300 14016 19306 14028
rect 19889 14025 19901 14028
rect 19935 14025 19947 14059
rect 19889 14019 19947 14025
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20901 14059 20959 14065
rect 20901 14056 20913 14059
rect 20680 14028 20913 14056
rect 20680 14016 20686 14028
rect 20901 14025 20913 14028
rect 20947 14025 20959 14059
rect 20901 14019 20959 14025
rect 12621 13991 12679 13997
rect 12621 13957 12633 13991
rect 12667 13957 12679 13991
rect 15010 13988 15016 14000
rect 12621 13951 12679 13957
rect 13280 13960 15016 13988
rect 13280 13932 13308 13960
rect 15010 13948 15016 13960
rect 15068 13948 15074 14000
rect 16390 13988 16396 14000
rect 16351 13960 16396 13988
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 17034 13948 17040 14000
rect 17092 13948 17098 14000
rect 17954 13948 17960 14000
rect 18012 13988 18018 14000
rect 18417 13991 18475 13997
rect 18417 13988 18429 13991
rect 18012 13960 18429 13988
rect 18012 13948 18018 13960
rect 18417 13957 18429 13960
rect 18463 13957 18475 13991
rect 18417 13951 18475 13957
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13920 8631 13923
rect 8662 13920 8668 13932
rect 8619 13892 8668 13920
rect 8619 13889 8631 13892
rect 8573 13883 8631 13889
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 13078 13920 13084 13932
rect 13039 13892 13084 13920
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13262 13920 13268 13932
rect 13223 13892 13268 13920
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13446 13920 13452 13932
rect 13407 13892 13452 13920
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13920 14151 13923
rect 14734 13920 14740 13932
rect 14139 13892 14740 13920
rect 14139 13889 14151 13892
rect 14093 13883 14151 13889
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 14826 13880 14832 13932
rect 14884 13920 14890 13932
rect 15102 13920 15108 13932
rect 14884 13892 14929 13920
rect 15063 13892 15108 13920
rect 14884 13880 14890 13892
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 16666 13920 16672 13932
rect 16627 13892 16672 13920
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 19058 13920 19064 13932
rect 19019 13892 19064 13920
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19208 13892 19441 13920
rect 19208 13880 19214 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19518 13880 19524 13932
rect 19576 13920 19582 13932
rect 20438 13920 20444 13932
rect 19576 13892 20444 13920
rect 19576 13880 19582 13892
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 14274 13852 14280 13864
rect 13955 13824 14280 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 14274 13812 14280 13824
rect 14332 13812 14338 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 15838 13852 15844 13864
rect 15611 13824 15844 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18877 13855 18935 13861
rect 18877 13852 18889 13855
rect 18196 13824 18889 13852
rect 18196 13812 18202 13824
rect 18877 13821 18889 13824
rect 18923 13821 18935 13855
rect 19334 13852 19340 13864
rect 19295 13824 19340 13852
rect 18877 13815 18935 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 8757 13787 8815 13793
rect 8757 13753 8769 13787
rect 8803 13784 8815 13787
rect 12710 13784 12716 13796
rect 8803 13756 12716 13784
rect 8803 13753 8815 13756
rect 8757 13747 8815 13753
rect 12710 13744 12716 13756
rect 12768 13784 12774 13796
rect 13446 13784 13452 13796
rect 12768 13756 13452 13784
rect 12768 13744 12774 13756
rect 13446 13744 13452 13756
rect 13504 13744 13510 13796
rect 13722 13744 13728 13796
rect 13780 13784 13786 13796
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 13780 13756 14933 13784
rect 13780 13744 13786 13756
rect 14921 13753 14933 13756
rect 14967 13784 14979 13787
rect 16574 13784 16580 13796
rect 14967 13756 16580 13784
rect 14967 13753 14979 13756
rect 14921 13747 14979 13753
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 20530 13744 20536 13796
rect 20588 13784 20594 13796
rect 20625 13787 20683 13793
rect 20625 13784 20637 13787
rect 20588 13756 20637 13784
rect 20588 13744 20594 13756
rect 20625 13753 20637 13756
rect 20671 13753 20683 13787
rect 20625 13747 20683 13753
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 15746 13676 15752 13728
rect 15804 13716 15810 13728
rect 15841 13719 15899 13725
rect 15841 13716 15853 13719
rect 15804 13688 15853 13716
rect 15804 13676 15810 13688
rect 15841 13685 15853 13688
rect 15887 13716 15899 13719
rect 15930 13716 15936 13728
rect 15887 13688 15936 13716
rect 15887 13685 15899 13688
rect 15841 13679 15899 13685
rect 15930 13676 15936 13688
rect 15988 13716 15994 13728
rect 17126 13716 17132 13728
rect 15988 13688 17132 13716
rect 15988 13676 15994 13688
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 21174 13676 21180 13728
rect 21232 13716 21238 13728
rect 21361 13719 21419 13725
rect 21361 13716 21373 13719
rect 21232 13688 21373 13716
rect 21232 13676 21238 13688
rect 21361 13685 21373 13688
rect 21407 13716 21419 13719
rect 21634 13716 21640 13728
rect 21407 13688 21640 13716
rect 21407 13685 21419 13688
rect 21361 13679 21419 13685
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 1104 13626 28336 13648
rect 1104 13574 3282 13626
rect 3334 13574 3346 13626
rect 3398 13574 3410 13626
rect 3462 13574 3474 13626
rect 3526 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 6410 13626
rect 6462 13574 6474 13626
rect 6526 13574 9282 13626
rect 9334 13574 9346 13626
rect 9398 13574 9410 13626
rect 9462 13574 9474 13626
rect 9526 13574 12282 13626
rect 12334 13574 12346 13626
rect 12398 13574 12410 13626
rect 12462 13574 12474 13626
rect 12526 13574 15282 13626
rect 15334 13574 15346 13626
rect 15398 13574 15410 13626
rect 15462 13574 15474 13626
rect 15526 13574 18282 13626
rect 18334 13574 18346 13626
rect 18398 13574 18410 13626
rect 18462 13574 18474 13626
rect 18526 13574 21282 13626
rect 21334 13574 21346 13626
rect 21398 13574 21410 13626
rect 21462 13574 21474 13626
rect 21526 13574 24282 13626
rect 24334 13574 24346 13626
rect 24398 13574 24410 13626
rect 24462 13574 24474 13626
rect 24526 13574 27282 13626
rect 27334 13574 27346 13626
rect 27398 13574 27410 13626
rect 27462 13574 27474 13626
rect 27526 13574 28336 13626
rect 1104 13552 28336 13574
rect 11977 13515 12035 13521
rect 11977 13481 11989 13515
rect 12023 13512 12035 13515
rect 12894 13512 12900 13524
rect 12023 13484 12900 13512
rect 12023 13481 12035 13484
rect 11977 13475 12035 13481
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 14826 13512 14832 13524
rect 14787 13484 14832 13512
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 15010 13472 15016 13524
rect 15068 13512 15074 13524
rect 15068 13484 15884 13512
rect 15068 13472 15074 13484
rect 10873 13447 10931 13453
rect 10873 13413 10885 13447
rect 10919 13444 10931 13447
rect 13262 13444 13268 13456
rect 10919 13416 13268 13444
rect 10919 13413 10931 13416
rect 10873 13407 10931 13413
rect 13262 13404 13268 13416
rect 13320 13404 13326 13456
rect 14553 13447 14611 13453
rect 14553 13413 14565 13447
rect 14599 13444 14611 13447
rect 15102 13444 15108 13456
rect 14599 13416 15108 13444
rect 14599 13413 14611 13416
rect 14553 13407 14611 13413
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 15749 13447 15807 13453
rect 15749 13413 15761 13447
rect 15795 13413 15807 13447
rect 15749 13407 15807 13413
rect 15856 13444 15884 13484
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 15988 13484 17325 13512
rect 15988 13472 15994 13484
rect 17313 13481 17325 13484
rect 17359 13481 17371 13515
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 17313 13475 17371 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 16853 13447 16911 13453
rect 16853 13444 16865 13447
rect 15856 13416 16865 13444
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13376 11667 13379
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 11655 13348 12909 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 12897 13345 12909 13348
rect 12943 13376 12955 13379
rect 13078 13376 13084 13388
rect 12943 13348 13084 13376
rect 12943 13345 12955 13348
rect 12897 13339 12955 13345
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 14182 13376 14188 13388
rect 13863 13348 14188 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 15620 13379 15678 13385
rect 15620 13376 15632 13379
rect 14976 13348 15632 13376
rect 14976 13336 14982 13348
rect 15620 13345 15632 13348
rect 15666 13345 15678 13379
rect 15620 13339 15678 13345
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 13357 13311 13415 13317
rect 11287 13280 13124 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 13096 13240 13124 13280
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13446 13308 13452 13320
rect 13403 13280 13452 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 13722 13308 13728 13320
rect 13683 13280 13728 13308
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 14274 13268 14280 13320
rect 14332 13308 14338 13320
rect 15764 13308 15792 13407
rect 15856 13385 15884 13416
rect 16853 13413 16865 13416
rect 16899 13444 16911 13447
rect 20898 13444 20904 13456
rect 16899 13416 20904 13444
rect 16899 13413 16911 13416
rect 16853 13407 16911 13413
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 16577 13379 16635 13385
rect 16577 13345 16589 13379
rect 16623 13376 16635 13379
rect 16666 13376 16672 13388
rect 16623 13348 16672 13376
rect 16623 13345 16635 13348
rect 16577 13339 16635 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 18877 13379 18935 13385
rect 18877 13345 18889 13379
rect 18923 13376 18935 13379
rect 19334 13376 19340 13388
rect 18923 13348 19340 13376
rect 18923 13345 18935 13348
rect 18877 13339 18935 13345
rect 19334 13336 19340 13348
rect 19392 13376 19398 13388
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 19392 13348 20085 13376
rect 19392 13336 19398 13348
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 17034 13308 17040 13320
rect 14332 13280 16436 13308
rect 16995 13280 17040 13308
rect 14332 13268 14338 13280
rect 14734 13240 14740 13252
rect 13096 13212 14740 13240
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 15473 13243 15531 13249
rect 15473 13209 15485 13243
rect 15519 13240 15531 13243
rect 15654 13240 15660 13252
rect 15519 13212 15660 13240
rect 15519 13209 15531 13212
rect 15473 13203 15531 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 16206 13240 16212 13252
rect 16167 13212 16212 13240
rect 16206 13200 16212 13212
rect 16264 13200 16270 13252
rect 16408 13240 16436 13280
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13308 17187 13311
rect 19058 13308 19064 13320
rect 17175 13280 18736 13308
rect 19019 13280 19064 13308
rect 17175 13277 17187 13280
rect 17129 13271 17187 13277
rect 17144 13240 17172 13271
rect 16408 13212 17172 13240
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 8573 13175 8631 13181
rect 8573 13172 8585 13175
rect 8444 13144 8585 13172
rect 8444 13132 8450 13144
rect 8573 13141 8585 13144
rect 8619 13172 8631 13175
rect 8662 13172 8668 13184
rect 8619 13144 8668 13172
rect 8619 13141 8631 13144
rect 8573 13135 8631 13141
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12710 13172 12716 13184
rect 12575 13144 12716 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 17957 13175 18015 13181
rect 17957 13141 17969 13175
rect 18003 13172 18015 13175
rect 18046 13172 18052 13184
rect 18003 13144 18052 13172
rect 18003 13141 18015 13144
rect 17957 13135 18015 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18138 13132 18144 13184
rect 18196 13172 18202 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 18196 13144 18245 13172
rect 18196 13132 18202 13144
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 18708 13172 18736 13280
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19150 13268 19156 13320
rect 19208 13308 19214 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 19208 13280 19257 13308
rect 19208 13268 19214 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 18874 13200 18880 13252
rect 18932 13240 18938 13252
rect 19628 13240 19656 13271
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 19760 13280 19805 13308
rect 19760 13268 19766 13280
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 22278 13308 22284 13320
rect 20404 13280 22284 13308
rect 20404 13268 20410 13280
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 22554 13240 22560 13252
rect 18932 13212 19656 13240
rect 22515 13212 22560 13240
rect 18932 13200 18938 13212
rect 22554 13200 22560 13212
rect 22612 13200 22618 13252
rect 23106 13200 23112 13252
rect 23164 13200 23170 13252
rect 23934 13200 23940 13252
rect 23992 13240 23998 13252
rect 24305 13243 24363 13249
rect 24305 13240 24317 13243
rect 23992 13212 24317 13240
rect 23992 13200 23998 13212
rect 24305 13209 24317 13212
rect 24351 13209 24363 13243
rect 24305 13203 24363 13209
rect 21085 13175 21143 13181
rect 21085 13172 21097 13175
rect 18708 13144 21097 13172
rect 18233 13135 18291 13141
rect 21085 13141 21097 13144
rect 21131 13141 21143 13175
rect 21085 13135 21143 13141
rect 21821 13175 21879 13181
rect 21821 13141 21833 13175
rect 21867 13172 21879 13175
rect 22462 13172 22468 13184
rect 21867 13144 22468 13172
rect 21867 13141 21879 13144
rect 21821 13135 21879 13141
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 1104 13082 28336 13104
rect 1104 13030 1782 13082
rect 1834 13030 1846 13082
rect 1898 13030 1910 13082
rect 1962 13030 1974 13082
rect 2026 13030 4782 13082
rect 4834 13030 4846 13082
rect 4898 13030 4910 13082
rect 4962 13030 4974 13082
rect 5026 13030 7782 13082
rect 7834 13030 7846 13082
rect 7898 13030 7910 13082
rect 7962 13030 7974 13082
rect 8026 13030 10782 13082
rect 10834 13030 10846 13082
rect 10898 13030 10910 13082
rect 10962 13030 10974 13082
rect 11026 13030 13782 13082
rect 13834 13030 13846 13082
rect 13898 13030 13910 13082
rect 13962 13030 13974 13082
rect 14026 13030 16782 13082
rect 16834 13030 16846 13082
rect 16898 13030 16910 13082
rect 16962 13030 16974 13082
rect 17026 13030 19782 13082
rect 19834 13030 19846 13082
rect 19898 13030 19910 13082
rect 19962 13030 19974 13082
rect 20026 13030 22782 13082
rect 22834 13030 22846 13082
rect 22898 13030 22910 13082
rect 22962 13030 22974 13082
rect 23026 13030 25782 13082
rect 25834 13030 25846 13082
rect 25898 13030 25910 13082
rect 25962 13030 25974 13082
rect 26026 13030 28336 13082
rect 1104 13008 28336 13030
rect 11238 12968 11244 12980
rect 11199 12940 11244 12968
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11701 12971 11759 12977
rect 11701 12937 11713 12971
rect 11747 12968 11759 12971
rect 13630 12968 13636 12980
rect 11747 12940 13636 12968
rect 11747 12937 11759 12940
rect 11701 12931 11759 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16482 12968 16488 12980
rect 16255 12940 16488 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 16945 12971 17003 12977
rect 16632 12940 16677 12968
rect 16632 12928 16638 12940
rect 16945 12937 16957 12971
rect 16991 12968 17003 12971
rect 17126 12968 17132 12980
rect 16991 12940 17132 12968
rect 16991 12937 17003 12940
rect 16945 12931 17003 12937
rect 14182 12900 14188 12912
rect 14095 12872 14188 12900
rect 14182 12860 14188 12872
rect 14240 12900 14246 12912
rect 16960 12900 16988 12931
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 19242 12968 19248 12980
rect 19203 12940 19248 12968
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21453 12971 21511 12977
rect 21453 12937 21465 12971
rect 21499 12968 21511 12971
rect 21726 12968 21732 12980
rect 21499 12940 21732 12968
rect 21499 12937 21511 12940
rect 21453 12931 21511 12937
rect 21726 12928 21732 12940
rect 21784 12968 21790 12980
rect 23106 12968 23112 12980
rect 21784 12940 23112 12968
rect 21784 12928 21790 12940
rect 23106 12928 23112 12940
rect 23164 12928 23170 12980
rect 23934 12968 23940 12980
rect 23895 12940 23940 12968
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 20162 12900 20168 12912
rect 14240 12872 16988 12900
rect 18892 12872 20168 12900
rect 14240 12860 14246 12872
rect 18892 12844 18920 12872
rect 20162 12860 20168 12872
rect 20220 12860 20226 12912
rect 22278 12860 22284 12912
rect 22336 12900 22342 12912
rect 23017 12903 23075 12909
rect 23017 12900 23029 12903
rect 22336 12872 23029 12900
rect 22336 12860 22342 12872
rect 23017 12869 23029 12872
rect 23063 12869 23075 12903
rect 23017 12863 23075 12869
rect 13262 12832 13268 12844
rect 13223 12804 13268 12832
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 13538 12832 13544 12844
rect 13499 12804 13544 12832
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15289 12835 15347 12841
rect 15289 12832 15301 12835
rect 15068 12804 15301 12832
rect 15068 12792 15074 12804
rect 15289 12801 15301 12804
rect 15335 12801 15347 12835
rect 15289 12795 15347 12801
rect 15657 12835 15715 12841
rect 15657 12801 15669 12835
rect 15703 12801 15715 12835
rect 15838 12832 15844 12844
rect 15799 12804 15844 12832
rect 15657 12795 15715 12801
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12115 12736 12909 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 13446 12764 13452 12776
rect 12943 12736 13452 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 14090 12764 14096 12776
rect 13863 12736 14096 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14700 12736 15209 12764
rect 14700 12724 14706 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 15672 12764 15700 12795
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 18782 12832 18788 12844
rect 18743 12804 18788 12832
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 18874 12792 18880 12844
rect 18932 12832 18938 12844
rect 18932 12804 18977 12832
rect 18932 12792 18938 12804
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 19334 12832 19340 12844
rect 19116 12804 19340 12832
rect 19116 12792 19122 12804
rect 19334 12792 19340 12804
rect 19392 12792 19398 12844
rect 22186 12832 22192 12844
rect 22147 12804 22192 12832
rect 22186 12792 22192 12804
rect 22244 12792 22250 12844
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 22520 12804 22569 12832
rect 22520 12792 22526 12804
rect 22557 12801 22569 12804
rect 22603 12832 22615 12835
rect 23952 12832 23980 12928
rect 22603 12804 23980 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 16482 12764 16488 12776
rect 15672 12736 16488 12764
rect 15197 12727 15255 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 18800 12764 18828 12792
rect 19150 12764 19156 12776
rect 18800 12736 19156 12764
rect 19150 12724 19156 12736
rect 19208 12764 19214 12776
rect 19797 12767 19855 12773
rect 19797 12764 19809 12767
rect 19208 12736 19809 12764
rect 19208 12724 19214 12736
rect 19797 12733 19809 12736
rect 19843 12733 19855 12767
rect 22646 12764 22652 12776
rect 22607 12736 22652 12764
rect 19797 12727 19855 12733
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 15562 12696 15568 12708
rect 13596 12668 15568 12696
rect 13596 12656 13602 12668
rect 15562 12656 15568 12668
rect 15620 12656 15626 12708
rect 18509 12699 18567 12705
rect 18509 12665 18521 12699
rect 18555 12696 18567 12699
rect 18690 12696 18696 12708
rect 18555 12668 18696 12696
rect 18555 12665 18567 12668
rect 18509 12659 18567 12665
rect 18690 12656 18696 12668
rect 18748 12696 18754 12708
rect 19610 12696 19616 12708
rect 18748 12668 19616 12696
rect 18748 12656 18754 12668
rect 19610 12656 19616 12668
rect 19668 12656 19674 12708
rect 22005 12699 22063 12705
rect 22005 12665 22017 12699
rect 22051 12696 22063 12699
rect 22554 12696 22560 12708
rect 22051 12668 22560 12696
rect 22051 12665 22063 12668
rect 22005 12659 22063 12665
rect 22554 12656 22560 12668
rect 22612 12656 22618 12708
rect 14737 12631 14795 12637
rect 14737 12597 14749 12631
rect 14783 12628 14795 12631
rect 15102 12628 15108 12640
rect 14783 12600 15108 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 17218 12628 17224 12640
rect 17179 12600 17224 12628
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17681 12631 17739 12637
rect 17681 12597 17693 12631
rect 17727 12628 17739 12631
rect 18046 12628 18052 12640
rect 17727 12600 18052 12628
rect 17727 12597 17739 12600
rect 17681 12591 17739 12597
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 20625 12631 20683 12637
rect 20625 12597 20637 12631
rect 20671 12628 20683 12631
rect 20714 12628 20720 12640
rect 20671 12600 20720 12628
rect 20671 12597 20683 12600
rect 20625 12591 20683 12597
rect 20714 12588 20720 12600
rect 20772 12628 20778 12640
rect 20990 12628 20996 12640
rect 20772 12600 20996 12628
rect 20772 12588 20778 12600
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 1104 12538 28336 12560
rect 1104 12486 3282 12538
rect 3334 12486 3346 12538
rect 3398 12486 3410 12538
rect 3462 12486 3474 12538
rect 3526 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 6410 12538
rect 6462 12486 6474 12538
rect 6526 12486 9282 12538
rect 9334 12486 9346 12538
rect 9398 12486 9410 12538
rect 9462 12486 9474 12538
rect 9526 12486 12282 12538
rect 12334 12486 12346 12538
rect 12398 12486 12410 12538
rect 12462 12486 12474 12538
rect 12526 12486 15282 12538
rect 15334 12486 15346 12538
rect 15398 12486 15410 12538
rect 15462 12486 15474 12538
rect 15526 12486 18282 12538
rect 18334 12486 18346 12538
rect 18398 12486 18410 12538
rect 18462 12486 18474 12538
rect 18526 12486 21282 12538
rect 21334 12486 21346 12538
rect 21398 12486 21410 12538
rect 21462 12486 21474 12538
rect 21526 12486 24282 12538
rect 24334 12486 24346 12538
rect 24398 12486 24410 12538
rect 24462 12486 24474 12538
rect 24526 12486 27282 12538
rect 27334 12486 27346 12538
rect 27398 12486 27410 12538
rect 27462 12486 27474 12538
rect 27526 12486 28336 12538
rect 1104 12464 28336 12486
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 13357 12427 13415 12433
rect 13357 12424 13369 12427
rect 8444 12396 13369 12424
rect 8444 12384 8450 12396
rect 13357 12393 13369 12396
rect 13403 12424 13415 12427
rect 13538 12424 13544 12436
rect 13403 12396 13544 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 15896 12396 17049 12424
rect 15896 12384 15902 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 17037 12387 17095 12393
rect 19613 12427 19671 12433
rect 19613 12393 19625 12427
rect 19659 12393 19671 12427
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 19613 12387 19671 12393
rect 15010 12316 15016 12368
rect 15068 12356 15074 12368
rect 15749 12359 15807 12365
rect 15749 12356 15761 12359
rect 15068 12328 15761 12356
rect 15068 12316 15074 12328
rect 15749 12325 15761 12328
rect 15795 12325 15807 12359
rect 15749 12319 15807 12325
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 19628 12356 19656 12387
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 22554 12424 22560 12436
rect 22515 12396 22560 12424
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 16724 12328 19656 12356
rect 16724 12316 16730 12328
rect 11054 12288 11060 12300
rect 10967 12260 11060 12288
rect 11054 12248 11060 12260
rect 11112 12288 11118 12300
rect 11882 12288 11888 12300
rect 11112 12260 11888 12288
rect 11112 12248 11118 12260
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 13228 12260 18337 12288
rect 13228 12248 13234 12260
rect 18325 12257 18337 12260
rect 18371 12257 18383 12291
rect 22186 12288 22192 12300
rect 22099 12260 22192 12288
rect 18325 12251 18383 12257
rect 22186 12248 22192 12260
rect 22244 12288 22250 12300
rect 22833 12291 22891 12297
rect 22833 12288 22845 12291
rect 22244 12260 22845 12288
rect 22244 12248 22250 12260
rect 22833 12257 22845 12260
rect 22879 12257 22891 12291
rect 23934 12288 23940 12300
rect 23895 12260 23940 12288
rect 22833 12251 22891 12257
rect 23934 12248 23940 12260
rect 23992 12248 23998 12300
rect 13262 12180 13268 12232
rect 13320 12220 13326 12232
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13320 12192 14197 12220
rect 13320 12180 13326 12192
rect 14185 12189 14197 12192
rect 14231 12220 14243 12223
rect 14458 12220 14464 12232
rect 14231 12192 14464 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14458 12180 14464 12192
rect 14516 12220 14522 12232
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 14516 12192 15485 12220
rect 14516 12180 14522 12192
rect 15473 12189 15485 12192
rect 15519 12220 15531 12223
rect 15930 12220 15936 12232
rect 15519 12192 15936 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 11330 12152 11336 12164
rect 11291 12124 11336 12152
rect 11330 12112 11336 12124
rect 11388 12112 11394 12164
rect 11790 12112 11796 12164
rect 11848 12112 11854 12164
rect 13081 12155 13139 12161
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 13538 12152 13544 12164
rect 13127 12124 13544 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 14274 12112 14280 12164
rect 14332 12152 14338 12164
rect 16408 12152 16436 12183
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 17586 12220 17592 12232
rect 16540 12192 16585 12220
rect 17547 12192 17592 12220
rect 16540 12180 16546 12192
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 18196 12192 18245 12220
rect 18196 12180 18202 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 19208 12192 19349 12220
rect 19208 12180 19214 12192
rect 19337 12189 19349 12192
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12220 19487 12223
rect 19518 12220 19524 12232
rect 19475 12192 19524 12220
rect 19475 12189 19487 12192
rect 19429 12183 19487 12189
rect 19518 12180 19524 12192
rect 19576 12180 19582 12232
rect 21726 12220 21732 12232
rect 21687 12192 21732 12220
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 17604 12152 17632 12180
rect 21928 12152 21956 12183
rect 22554 12152 22560 12164
rect 14332 12124 17632 12152
rect 21100 12124 22560 12152
rect 14332 12112 14338 12124
rect 21100 12096 21128 12124
rect 22554 12112 22560 12124
rect 22612 12112 22618 12164
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10652 12056 10701 12084
rect 10652 12044 10658 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13504 12056 13829 12084
rect 13504 12044 13510 12056
rect 13817 12053 13829 12056
rect 13863 12084 13875 12087
rect 14642 12084 14648 12096
rect 13863 12056 14648 12084
rect 13863 12053 13875 12056
rect 13817 12047 13875 12053
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 18782 12044 18788 12096
rect 18840 12084 18846 12096
rect 18877 12087 18935 12093
rect 18877 12084 18889 12087
rect 18840 12056 18889 12084
rect 18840 12044 18846 12056
rect 18877 12053 18889 12056
rect 18923 12084 18935 12087
rect 19058 12084 19064 12096
rect 18923 12056 19064 12084
rect 18923 12053 18935 12056
rect 18877 12047 18935 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 21082 12084 21088 12096
rect 21043 12056 21088 12084
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 23474 12044 23480 12096
rect 23532 12084 23538 12096
rect 24302 12084 24308 12096
rect 23532 12056 24308 12084
rect 23532 12044 23538 12056
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 1104 11994 28336 12016
rect 1104 11942 1782 11994
rect 1834 11942 1846 11994
rect 1898 11942 1910 11994
rect 1962 11942 1974 11994
rect 2026 11942 4782 11994
rect 4834 11942 4846 11994
rect 4898 11942 4910 11994
rect 4962 11942 4974 11994
rect 5026 11942 7782 11994
rect 7834 11942 7846 11994
rect 7898 11942 7910 11994
rect 7962 11942 7974 11994
rect 8026 11942 10782 11994
rect 10834 11942 10846 11994
rect 10898 11942 10910 11994
rect 10962 11942 10974 11994
rect 11026 11942 13782 11994
rect 13834 11942 13846 11994
rect 13898 11942 13910 11994
rect 13962 11942 13974 11994
rect 14026 11942 16782 11994
rect 16834 11942 16846 11994
rect 16898 11942 16910 11994
rect 16962 11942 16974 11994
rect 17026 11942 19782 11994
rect 19834 11942 19846 11994
rect 19898 11942 19910 11994
rect 19962 11942 19974 11994
rect 20026 11942 22782 11994
rect 22834 11942 22846 11994
rect 22898 11942 22910 11994
rect 22962 11942 22974 11994
rect 23026 11960 25782 11994
rect 23026 11942 24308 11960
rect 1104 11920 24308 11942
rect 24302 11908 24308 11920
rect 24360 11942 25782 11960
rect 25834 11942 25846 11994
rect 25898 11942 25910 11994
rect 25962 11942 25974 11994
rect 26026 11942 28336 11994
rect 24360 11920 28336 11942
rect 24360 11908 24366 11920
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 10652 11852 10701 11880
rect 10652 11840 10658 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 11146 11880 11152 11892
rect 11107 11852 11152 11880
rect 10689 11843 10747 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 11388 11852 11437 11880
rect 11388 11840 11394 11852
rect 11425 11849 11437 11852
rect 11471 11880 11483 11883
rect 14458 11880 14464 11892
rect 11471 11852 12664 11880
rect 14419 11852 14464 11880
rect 11471 11849 11483 11852
rect 11425 11843 11483 11849
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 11164 11812 11192 11840
rect 11790 11812 11796 11824
rect 10468 11784 11192 11812
rect 11751 11784 11796 11812
rect 10468 11772 10474 11784
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 12636 11821 12664 11852
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 16080 11852 17049 11880
rect 16080 11840 16086 11852
rect 17037 11849 17049 11852
rect 17083 11880 17095 11883
rect 17083 11852 17540 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 12621 11815 12679 11821
rect 12621 11781 12633 11815
rect 12667 11781 12679 11815
rect 14182 11812 14188 11824
rect 12621 11775 12679 11781
rect 13280 11784 14188 11812
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8938 11744 8944 11756
rect 8159 11716 8944 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 13170 11744 13176 11756
rect 13131 11716 13176 11744
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 13280 11753 13308 11784
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 15654 11812 15660 11824
rect 15488 11784 15660 11812
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11713 13323 11747
rect 13446 11744 13452 11756
rect 13407 11716 13452 11744
rect 13265 11707 13323 11713
rect 8018 11676 8024 11688
rect 7979 11648 8024 11676
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 12618 11676 12624 11688
rect 11296 11648 12624 11676
rect 11296 11636 11302 11648
rect 12618 11636 12624 11648
rect 12676 11676 12682 11688
rect 13280 11676 13308 11707
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 14090 11744 14096 11756
rect 14051 11716 14096 11744
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15488 11753 15516 11784
rect 15654 11772 15660 11784
rect 15712 11812 15718 11824
rect 17218 11812 17224 11824
rect 15712 11784 17224 11812
rect 15712 11772 15718 11784
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 17512 11812 17540 11852
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 22554 11880 22560 11892
rect 17644 11852 19656 11880
rect 22515 11852 22560 11880
rect 17644 11840 17650 11852
rect 17770 11812 17776 11824
rect 17512 11784 17776 11812
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 19628 11812 19656 11852
rect 22554 11840 22560 11852
rect 22612 11840 22618 11892
rect 22925 11815 22983 11821
rect 22925 11812 22937 11815
rect 19628 11784 22937 11812
rect 22925 11781 22937 11784
rect 22971 11781 22983 11815
rect 22925 11775 22983 11781
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 15160 11716 15209 11744
rect 15160 11704 15166 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 18690 11744 18696 11756
rect 15620 11716 15665 11744
rect 18651 11716 18696 11744
rect 15620 11704 15626 11716
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 18923 11716 19104 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 12676 11648 13308 11676
rect 12676 11636 12682 11648
rect 13538 11636 13544 11688
rect 13596 11676 13602 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13596 11648 13921 11676
rect 13596 11636 13602 11648
rect 13909 11645 13921 11648
rect 13955 11676 13967 11679
rect 14274 11676 14280 11688
rect 13955 11648 14280 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14734 11676 14740 11688
rect 14695 11648 14740 11676
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15488 11648 15853 11676
rect 13722 11568 13728 11620
rect 13780 11608 13786 11620
rect 15488 11608 15516 11648
rect 15841 11645 15853 11648
rect 15887 11645 15899 11679
rect 16114 11676 16120 11688
rect 16075 11648 16120 11676
rect 15841 11639 15899 11645
rect 16114 11636 16120 11648
rect 16172 11676 16178 11688
rect 16482 11676 16488 11688
rect 16172 11648 16488 11676
rect 16172 11636 16178 11648
rect 16482 11636 16488 11648
rect 16540 11676 16546 11688
rect 17126 11676 17132 11688
rect 16540 11648 17132 11676
rect 16540 11636 16546 11648
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18414 11676 18420 11688
rect 18104 11648 18420 11676
rect 18104 11636 18110 11648
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 13780 11580 15516 11608
rect 13780 11568 13786 11580
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 8297 11543 8355 11549
rect 8297 11540 8309 11543
rect 6236 11512 8309 11540
rect 6236 11500 6242 11512
rect 8297 11509 8309 11512
rect 8343 11509 8355 11543
rect 8297 11503 8355 11509
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 14976 11512 16497 11540
rect 14976 11500 14982 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 17494 11540 17500 11552
rect 17455 11512 17500 11540
rect 16485 11503 16543 11509
rect 17494 11500 17500 11512
rect 17552 11540 17558 11552
rect 18138 11540 18144 11552
rect 17552 11512 18144 11540
rect 17552 11500 17558 11512
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 19076 11540 19104 11716
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19337 11747 19395 11753
rect 19337 11744 19349 11747
rect 19300 11716 19349 11744
rect 19300 11704 19306 11716
rect 19337 11713 19349 11716
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 21726 11744 21732 11756
rect 19484 11716 21496 11744
rect 21639 11716 21732 11744
rect 19484 11704 19490 11716
rect 20898 11676 20904 11688
rect 20859 11648 20904 11676
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 21468 11685 21496 11716
rect 21726 11704 21732 11716
rect 21784 11744 21790 11756
rect 22278 11744 22284 11756
rect 21784 11716 22284 11744
rect 21784 11704 21790 11716
rect 22278 11704 22284 11716
rect 22336 11704 22342 11756
rect 21453 11679 21511 11685
rect 21453 11645 21465 11679
rect 21499 11676 21511 11679
rect 21818 11676 21824 11688
rect 21499 11648 21824 11676
rect 21499 11645 21511 11648
rect 21453 11639 21511 11645
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 21913 11679 21971 11685
rect 21913 11645 21925 11679
rect 21959 11645 21971 11679
rect 21913 11639 21971 11645
rect 25041 11679 25099 11685
rect 25041 11645 25053 11679
rect 25087 11676 25099 11679
rect 28718 11676 28724 11688
rect 25087 11648 28724 11676
rect 25087 11645 25099 11648
rect 25041 11639 25099 11645
rect 19794 11608 19800 11620
rect 19755 11580 19800 11608
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 20990 11608 20996 11620
rect 20272 11580 20996 11608
rect 20272 11540 20300 11580
rect 20990 11568 20996 11580
rect 21048 11568 21054 11620
rect 19076 11512 20300 11540
rect 20346 11500 20352 11552
rect 20404 11540 20410 11552
rect 21928 11540 21956 11639
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 22278 11540 22284 11552
rect 20404 11512 21956 11540
rect 22239 11512 22284 11540
rect 20404 11500 20410 11512
rect 22278 11500 22284 11512
rect 22336 11500 22342 11552
rect 1104 11450 28336 11472
rect 1104 11398 3282 11450
rect 3334 11398 3346 11450
rect 3398 11398 3410 11450
rect 3462 11398 3474 11450
rect 3526 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 6410 11450
rect 6462 11398 6474 11450
rect 6526 11398 9282 11450
rect 9334 11398 9346 11450
rect 9398 11398 9410 11450
rect 9462 11398 9474 11450
rect 9526 11398 12282 11450
rect 12334 11398 12346 11450
rect 12398 11398 12410 11450
rect 12462 11398 12474 11450
rect 12526 11398 15282 11450
rect 15334 11398 15346 11450
rect 15398 11398 15410 11450
rect 15462 11398 15474 11450
rect 15526 11398 18282 11450
rect 18334 11398 18346 11450
rect 18398 11398 18410 11450
rect 18462 11398 18474 11450
rect 18526 11398 21282 11450
rect 21334 11398 21346 11450
rect 21398 11398 21410 11450
rect 21462 11398 21474 11450
rect 21526 11398 24282 11450
rect 24334 11398 24346 11450
rect 24398 11398 24410 11450
rect 24462 11398 24474 11450
rect 24526 11398 27282 11450
rect 27334 11398 27346 11450
rect 27398 11398 27410 11450
rect 27462 11398 27474 11450
rect 27526 11398 28336 11450
rect 1104 11376 28336 11398
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 11790 11336 11796 11348
rect 11103 11308 11796 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11336 12955 11339
rect 13170 11336 13176 11348
rect 12943 11308 13176 11336
rect 12943 11305 12955 11308
rect 12897 11299 12955 11305
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 14090 11336 14096 11348
rect 13311 11308 14096 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 15102 11296 15108 11348
rect 15160 11336 15166 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15160 11308 15945 11336
rect 15160 11296 15166 11308
rect 15933 11305 15945 11308
rect 15979 11305 15991 11339
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 15933 11299 15991 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18417 11339 18475 11345
rect 18417 11305 18429 11339
rect 18463 11336 18475 11339
rect 19242 11336 19248 11348
rect 18463 11308 19248 11336
rect 18463 11305 18475 11308
rect 18417 11299 18475 11305
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19518 11336 19524 11348
rect 19431 11308 19524 11336
rect 19518 11296 19524 11308
rect 19576 11336 19582 11348
rect 19794 11336 19800 11348
rect 19576 11308 19800 11336
rect 19576 11296 19582 11308
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 21082 11336 21088 11348
rect 19935 11308 21088 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 12069 11271 12127 11277
rect 12069 11237 12081 11271
rect 12115 11268 12127 11271
rect 13722 11268 13728 11280
rect 12115 11240 13728 11268
rect 12115 11237 12127 11240
rect 12069 11231 12127 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 14461 11271 14519 11277
rect 14461 11237 14473 11271
rect 14507 11268 14519 11271
rect 15654 11268 15660 11280
rect 14507 11240 15660 11268
rect 14507 11237 14519 11240
rect 14461 11231 14519 11237
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 16761 11271 16819 11277
rect 16761 11237 16773 11271
rect 16807 11268 16819 11271
rect 17218 11268 17224 11280
rect 16807 11240 17224 11268
rect 16807 11237 16819 11240
rect 16761 11231 16819 11237
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 18782 11268 18788 11280
rect 18743 11240 18788 11268
rect 18782 11228 18788 11240
rect 18840 11228 18846 11280
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 12437 11203 12495 11209
rect 12437 11200 12449 11203
rect 11388 11172 12449 11200
rect 11388 11160 11394 11172
rect 12437 11169 12449 11172
rect 12483 11200 12495 11203
rect 12710 11200 12716 11212
rect 12483 11172 12716 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 12710 11160 12716 11172
rect 12768 11200 12774 11212
rect 13446 11200 13452 11212
rect 12768 11172 13452 11200
rect 12768 11160 12774 11172
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 14093 11203 14151 11209
rect 14093 11169 14105 11203
rect 14139 11200 14151 11203
rect 15010 11200 15016 11212
rect 14139 11172 15016 11200
rect 14139 11169 14151 11172
rect 14093 11163 14151 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 17586 11200 17592 11212
rect 16960 11172 17592 11200
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9030 11132 9036 11144
rect 8803 11104 9036 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 7745 11067 7803 11073
rect 7745 11033 7757 11067
rect 7791 11064 7803 11067
rect 8018 11064 8024 11076
rect 7791 11036 8024 11064
rect 7791 11033 7803 11036
rect 7745 11027 7803 11033
rect 8018 11024 8024 11036
rect 8076 11064 8082 11076
rect 8772 11064 8800 11095
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11146 11132 11152 11144
rect 10919 11104 11152 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 11974 11132 11980 11144
rect 11931 11104 11980 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 11974 11092 11980 11104
rect 12032 11092 12038 11144
rect 15470 11132 15476 11144
rect 15431 11104 15476 11132
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 16960 11141 16988 11172
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 19610 11200 19616 11212
rect 19571 11172 19616 11200
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 21818 11200 21824 11212
rect 21731 11172 21824 11200
rect 21818 11160 21824 11172
rect 21876 11200 21882 11212
rect 22097 11203 22155 11209
rect 22097 11200 22109 11203
rect 21876 11172 22109 11200
rect 21876 11160 21882 11172
rect 22097 11169 22109 11172
rect 22143 11169 22155 11203
rect 22097 11163 22155 11169
rect 22278 11160 22284 11212
rect 22336 11200 22342 11212
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 22336 11172 22477 11200
rect 22336 11160 22342 11172
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 22465 11163 22523 11169
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11101 17003 11135
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 16945 11095 17003 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17678 11092 17684 11144
rect 17736 11132 17742 11144
rect 19392 11135 19450 11141
rect 19392 11132 19404 11135
rect 17736 11104 19404 11132
rect 17736 11092 17742 11104
rect 19392 11101 19404 11104
rect 19438 11132 19450 11135
rect 20898 11132 20904 11144
rect 19438 11104 20904 11132
rect 19438 11101 19450 11104
rect 19392 11095 19450 11101
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 21726 11132 21732 11144
rect 21687 11104 21732 11132
rect 21726 11092 21732 11104
rect 21784 11092 21790 11144
rect 22557 11135 22615 11141
rect 22557 11101 22569 11135
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 8076 11036 8800 11064
rect 14829 11067 14887 11073
rect 8076 11024 8082 11036
rect 14829 11033 14841 11067
rect 14875 11064 14887 11067
rect 15562 11064 15568 11076
rect 14875 11036 15568 11064
rect 14875 11033 14887 11036
rect 14829 11027 14887 11033
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 16264 11036 19257 11064
rect 16264 11024 16270 11036
rect 19245 11033 19257 11036
rect 19291 11064 19303 11067
rect 21174 11064 21180 11076
rect 19291 11036 21180 11064
rect 19291 11033 19303 11036
rect 19245 11027 19303 11033
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 22462 11024 22468 11076
rect 22520 11064 22526 11076
rect 22572 11064 22600 11095
rect 22520 11036 22600 11064
rect 22520 11024 22526 11036
rect 6914 10996 6920 11008
rect 6875 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 8938 10956 8944 11008
rect 8996 10996 9002 11008
rect 9033 10999 9091 11005
rect 9033 10996 9045 10999
rect 8996 10968 9045 10996
rect 8996 10956 9002 10968
rect 9033 10965 9045 10968
rect 9079 10965 9091 10999
rect 11606 10996 11612 11008
rect 11567 10968 11612 10996
rect 9033 10959 9091 10965
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 15657 10999 15715 11005
rect 15657 10965 15669 10999
rect 15703 10996 15715 10999
rect 19150 10996 19156 11008
rect 15703 10968 19156 10996
rect 15703 10965 15715 10968
rect 15657 10959 15715 10965
rect 19150 10956 19156 10968
rect 19208 10996 19214 11008
rect 20346 10996 20352 11008
rect 19208 10968 20352 10996
rect 19208 10956 19214 10968
rect 20346 10956 20352 10968
rect 20404 10996 20410 11008
rect 20441 10999 20499 11005
rect 20441 10996 20453 10999
rect 20404 10968 20453 10996
rect 20404 10956 20410 10968
rect 20441 10965 20453 10968
rect 20487 10965 20499 10999
rect 20441 10959 20499 10965
rect 1104 10906 28336 10928
rect 1104 10854 1782 10906
rect 1834 10854 1846 10906
rect 1898 10854 1910 10906
rect 1962 10854 1974 10906
rect 2026 10854 4782 10906
rect 4834 10854 4846 10906
rect 4898 10854 4910 10906
rect 4962 10854 4974 10906
rect 5026 10854 7782 10906
rect 7834 10854 7846 10906
rect 7898 10854 7910 10906
rect 7962 10854 7974 10906
rect 8026 10854 10782 10906
rect 10834 10854 10846 10906
rect 10898 10854 10910 10906
rect 10962 10854 10974 10906
rect 11026 10854 13782 10906
rect 13834 10854 13846 10906
rect 13898 10854 13910 10906
rect 13962 10854 13974 10906
rect 14026 10854 16782 10906
rect 16834 10854 16846 10906
rect 16898 10854 16910 10906
rect 16962 10854 16974 10906
rect 17026 10854 19782 10906
rect 19834 10854 19846 10906
rect 19898 10854 19910 10906
rect 19962 10854 19974 10906
rect 20026 10854 22782 10906
rect 22834 10854 22846 10906
rect 22898 10854 22910 10906
rect 22962 10854 22974 10906
rect 23026 10854 25782 10906
rect 25834 10854 25846 10906
rect 25898 10854 25910 10906
rect 25962 10854 25974 10906
rect 26026 10854 28336 10906
rect 1104 10832 28336 10854
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 8110 10792 8116 10804
rect 6503 10764 8116 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11146 10792 11152 10804
rect 11103 10764 11152 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 13081 10795 13139 10801
rect 13081 10792 13093 10795
rect 11664 10764 13093 10792
rect 11664 10752 11670 10764
rect 13081 10761 13093 10764
rect 13127 10792 13139 10795
rect 13449 10795 13507 10801
rect 13449 10792 13461 10795
rect 13127 10764 13461 10792
rect 13127 10761 13139 10764
rect 13081 10755 13139 10761
rect 13449 10761 13461 10764
rect 13495 10792 13507 10795
rect 13538 10792 13544 10804
rect 13495 10764 13544 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 17678 10792 17684 10804
rect 17639 10764 17684 10792
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 17770 10752 17776 10804
rect 17828 10792 17834 10804
rect 19426 10792 19432 10804
rect 17828 10764 19432 10792
rect 17828 10752 17834 10764
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 19610 10752 19616 10804
rect 19668 10792 19674 10804
rect 19705 10795 19763 10801
rect 19705 10792 19717 10795
rect 19668 10764 19717 10792
rect 19668 10752 19674 10764
rect 19705 10761 19717 10764
rect 19751 10792 19763 10795
rect 21821 10795 21879 10801
rect 19751 10764 20300 10792
rect 19751 10761 19763 10764
rect 19705 10755 19763 10761
rect 12618 10724 12624 10736
rect 12579 10696 12624 10724
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 14550 10684 14556 10736
rect 14608 10684 14614 10736
rect 15470 10684 15476 10736
rect 15528 10724 15534 10736
rect 16209 10727 16267 10733
rect 16209 10724 16221 10727
rect 15528 10696 16221 10724
rect 15528 10684 15534 10696
rect 16209 10693 16221 10696
rect 16255 10724 16267 10727
rect 17310 10724 17316 10736
rect 16255 10696 17316 10724
rect 16255 10693 16267 10696
rect 16209 10687 16267 10693
rect 17310 10684 17316 10696
rect 17368 10724 17374 10736
rect 18969 10727 19027 10733
rect 18969 10724 18981 10727
rect 17368 10696 18981 10724
rect 17368 10684 17374 10696
rect 18969 10693 18981 10696
rect 19015 10724 19027 10727
rect 19242 10724 19248 10736
rect 19015 10696 19248 10724
rect 19015 10693 19027 10696
rect 18969 10687 19027 10693
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 20272 10733 20300 10764
rect 21821 10761 21833 10795
rect 21867 10792 21879 10795
rect 22278 10792 22284 10804
rect 21867 10764 22284 10792
rect 21867 10761 21879 10764
rect 21821 10755 21879 10761
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 20257 10727 20315 10733
rect 20257 10693 20269 10727
rect 20303 10693 20315 10727
rect 20257 10687 20315 10693
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 7484 10628 8401 10656
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7484 10461 7512 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8938 10656 8944 10668
rect 8389 10619 8447 10625
rect 8496 10628 8944 10656
rect 8294 10588 8300 10600
rect 8255 10560 8300 10588
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8496 10520 8524 10628
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 9088 10628 9137 10656
rect 9088 10616 9094 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 10376 10628 10517 10656
rect 10376 10616 10382 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 13538 10656 13544 10668
rect 11940 10628 13544 10656
rect 11940 10616 11946 10628
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 16761 10659 16819 10665
rect 13596 10628 13860 10656
rect 13596 10616 13602 10628
rect 13832 10597 13860 10628
rect 16761 10625 16773 10659
rect 16807 10625 16819 10659
rect 18874 10656 18880 10668
rect 18835 10628 18880 10656
rect 16761 10619 16819 10625
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 14734 10588 14740 10600
rect 14139 10560 14740 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 15841 10591 15899 10597
rect 15841 10557 15853 10591
rect 15887 10588 15899 10591
rect 16206 10588 16212 10600
rect 15887 10560 16212 10588
rect 15887 10557 15899 10560
rect 15841 10551 15899 10557
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16776 10588 16804 10619
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 20898 10656 20904 10668
rect 20859 10628 20904 10656
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 21726 10656 21732 10668
rect 21315 10628 21732 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21726 10616 21732 10628
rect 21784 10656 21790 10668
rect 21784 10628 22232 10656
rect 21784 10616 21790 10628
rect 18966 10588 18972 10600
rect 16356 10560 18972 10588
rect 16356 10548 16362 10560
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 20070 10548 20076 10600
rect 20128 10588 20134 10600
rect 20809 10591 20867 10597
rect 20809 10588 20821 10591
rect 20128 10560 20821 10588
rect 20128 10548 20134 10560
rect 20809 10557 20821 10560
rect 20855 10557 20867 10591
rect 20809 10551 20867 10557
rect 20990 10548 20996 10600
rect 21048 10588 21054 10600
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 21048 10560 21373 10588
rect 21048 10548 21054 10560
rect 21361 10557 21373 10560
rect 21407 10588 21419 10591
rect 21910 10588 21916 10600
rect 21407 10560 21916 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 7852 10492 8524 10520
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6788 10424 7021 10452
rect 6788 10412 6794 10424
rect 7009 10421 7021 10424
rect 7055 10452 7067 10455
rect 7469 10455 7527 10461
rect 7469 10452 7481 10455
rect 7055 10424 7481 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7469 10421 7481 10424
rect 7515 10421 7527 10455
rect 7469 10415 7527 10421
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7852 10461 7880 10492
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 9309 10523 9367 10529
rect 9309 10520 9321 10523
rect 9180 10492 9321 10520
rect 9180 10480 9186 10492
rect 9309 10489 9321 10492
rect 9355 10489 9367 10523
rect 9309 10483 9367 10489
rect 10689 10523 10747 10529
rect 10689 10489 10701 10523
rect 10735 10520 10747 10523
rect 11146 10520 11152 10532
rect 10735 10492 11152 10520
rect 10735 10489 10747 10492
rect 10689 10483 10747 10489
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 22204 10520 22232 10628
rect 22833 10523 22891 10529
rect 22833 10520 22845 10523
rect 22204 10492 22845 10520
rect 22204 10464 22232 10492
rect 22833 10489 22845 10492
rect 22879 10520 22891 10523
rect 23842 10520 23848 10532
rect 22879 10492 23848 10520
rect 22879 10489 22891 10492
rect 22833 10483 22891 10489
rect 23842 10480 23848 10492
rect 23900 10480 23906 10532
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7708 10424 7849 10452
rect 7708 10412 7714 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 7837 10415 7895 10421
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9582 10452 9588 10464
rect 8352 10424 9588 10452
rect 8352 10412 8358 10424
rect 9582 10412 9588 10424
rect 9640 10452 9646 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 9640 10424 9873 10452
rect 9640 10412 9646 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 11974 10452 11980 10464
rect 11935 10424 11980 10452
rect 9861 10415 9919 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 13814 10452 13820 10464
rect 13044 10424 13820 10452
rect 13044 10412 13050 10424
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 15838 10412 15844 10464
rect 15896 10452 15902 10464
rect 16945 10455 17003 10461
rect 16945 10452 16957 10455
rect 15896 10424 16957 10452
rect 15896 10412 15902 10424
rect 16945 10421 16957 10424
rect 16991 10452 17003 10455
rect 21634 10452 21640 10464
rect 16991 10424 21640 10452
rect 16991 10421 17003 10424
rect 16945 10415 17003 10421
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 22186 10452 22192 10464
rect 22147 10424 22192 10452
rect 22186 10412 22192 10424
rect 22244 10412 22250 10464
rect 22462 10452 22468 10464
rect 22423 10424 22468 10452
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 1104 10362 28336 10384
rect 1104 10310 3282 10362
rect 3334 10310 3346 10362
rect 3398 10310 3410 10362
rect 3462 10310 3474 10362
rect 3526 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 6410 10362
rect 6462 10310 6474 10362
rect 6526 10310 9282 10362
rect 9334 10310 9346 10362
rect 9398 10310 9410 10362
rect 9462 10310 9474 10362
rect 9526 10310 12282 10362
rect 12334 10310 12346 10362
rect 12398 10310 12410 10362
rect 12462 10310 12474 10362
rect 12526 10310 15282 10362
rect 15334 10310 15346 10362
rect 15398 10310 15410 10362
rect 15462 10310 15474 10362
rect 15526 10310 18282 10362
rect 18334 10310 18346 10362
rect 18398 10310 18410 10362
rect 18462 10310 18474 10362
rect 18526 10310 21282 10362
rect 21334 10310 21346 10362
rect 21398 10310 21410 10362
rect 21462 10310 21474 10362
rect 21526 10310 24282 10362
rect 24334 10310 24346 10362
rect 24398 10310 24410 10362
rect 24462 10310 24474 10362
rect 24526 10310 27282 10362
rect 27334 10310 27346 10362
rect 27398 10310 27410 10362
rect 27462 10310 27474 10362
rect 27526 10310 28336 10362
rect 1104 10288 28336 10310
rect 6365 10251 6423 10257
rect 6365 10217 6377 10251
rect 6411 10248 6423 10251
rect 6730 10248 6736 10260
rect 6411 10220 6736 10248
rect 6411 10217 6423 10220
rect 6365 10211 6423 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 6914 10248 6920 10260
rect 6875 10220 6920 10248
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 9030 10248 9036 10260
rect 8991 10220 9036 10248
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 12986 10248 12992 10260
rect 10744 10220 12992 10248
rect 10744 10208 10750 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10248 13507 10251
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 13495 10220 13921 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 13909 10217 13921 10220
rect 13955 10248 13967 10251
rect 14550 10248 14556 10260
rect 13955 10220 14556 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 14645 10251 14703 10257
rect 14645 10217 14657 10251
rect 14691 10248 14703 10251
rect 14734 10248 14740 10260
rect 14691 10220 14740 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14884 10220 16436 10248
rect 14884 10208 14890 10220
rect 8294 10180 8300 10192
rect 8220 10152 8300 10180
rect 8220 10112 8248 10152
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12032 10152 16344 10180
rect 12032 10140 12038 10152
rect 10410 10112 10416 10124
rect 7944 10084 8248 10112
rect 10371 10084 10416 10112
rect 6178 10044 6184 10056
rect 6139 10016 6184 10044
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6914 10004 6920 10056
rect 6972 10044 6978 10056
rect 7944 10053 7972 10084
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 16206 10112 16212 10124
rect 13872 10084 16212 10112
rect 13872 10072 13878 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 6972 10016 7665 10044
rect 6972 10004 6978 10016
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8294 10044 8300 10056
rect 8255 10016 8300 10044
rect 8021 10007 8079 10013
rect 7193 9979 7251 9985
rect 7193 9945 7205 9979
rect 7239 9976 7251 9979
rect 7282 9976 7288 9988
rect 7239 9948 7288 9976
rect 7239 9945 7251 9948
rect 7193 9939 7251 9945
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 7558 9936 7564 9988
rect 7616 9976 7622 9988
rect 8036 9976 8064 10007
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13412 10016 13737 10044
rect 13412 10004 13418 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 15654 10044 15660 10056
rect 15615 10016 15660 10044
rect 13725 10007 13783 10013
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 16316 10044 16344 10152
rect 16408 10112 16436 10220
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 16724 10220 17509 10248
rect 16724 10208 16730 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 17497 10211 17555 10217
rect 18049 10251 18107 10257
rect 18049 10217 18061 10251
rect 18095 10248 18107 10251
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 18095 10220 18981 10248
rect 18095 10217 18107 10220
rect 18049 10211 18107 10217
rect 18969 10217 18981 10220
rect 19015 10217 19027 10251
rect 18969 10211 19027 10217
rect 18984 10180 19012 10211
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19576 10220 19717 10248
rect 19576 10208 19582 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 19705 10211 19763 10217
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21453 10251 21511 10257
rect 21453 10248 21465 10251
rect 21232 10220 21465 10248
rect 21232 10208 21238 10220
rect 21453 10217 21465 10220
rect 21499 10217 21511 10251
rect 21453 10211 21511 10217
rect 20530 10180 20536 10192
rect 18984 10152 20536 10180
rect 20530 10140 20536 10152
rect 20588 10180 20594 10192
rect 20898 10180 20904 10192
rect 20588 10152 20904 10180
rect 20588 10140 20594 10152
rect 20898 10140 20904 10152
rect 20956 10180 20962 10192
rect 21085 10183 21143 10189
rect 21085 10180 21097 10183
rect 20956 10152 21097 10180
rect 20956 10140 20962 10152
rect 21085 10149 21097 10152
rect 21131 10149 21143 10183
rect 21085 10143 21143 10149
rect 17129 10115 17187 10121
rect 17129 10112 17141 10115
rect 16408 10084 17141 10112
rect 17129 10081 17141 10084
rect 17175 10081 17187 10115
rect 17129 10075 17187 10081
rect 19061 10115 19119 10121
rect 19061 10081 19073 10115
rect 19107 10112 19119 10115
rect 20070 10112 20076 10124
rect 19107 10084 20076 10112
rect 19107 10081 19119 10084
rect 19061 10075 19119 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21821 10115 21879 10121
rect 21821 10112 21833 10115
rect 20772 10084 21833 10112
rect 20772 10072 20778 10084
rect 21821 10081 21833 10084
rect 21867 10112 21879 10115
rect 22094 10112 22100 10124
rect 21867 10084 22100 10112
rect 21867 10081 21879 10084
rect 21821 10075 21879 10081
rect 22094 10072 22100 10084
rect 22152 10072 22158 10124
rect 23842 10112 23848 10124
rect 23803 10084 23848 10112
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 16393 10047 16451 10053
rect 16393 10044 16405 10047
rect 16316 10016 16405 10044
rect 16393 10013 16405 10016
rect 16439 10044 16451 10047
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16439 10016 16865 10044
rect 16439 10013 16451 10016
rect 16393 10007 16451 10013
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 18417 10047 18475 10053
rect 18417 10013 18429 10047
rect 18463 10044 18475 10047
rect 18840 10047 18898 10053
rect 18840 10044 18852 10047
rect 18463 10016 18852 10044
rect 18463 10013 18475 10016
rect 18417 10007 18475 10013
rect 18840 10013 18852 10016
rect 18886 10044 18898 10047
rect 19518 10044 19524 10056
rect 18886 10016 19524 10044
rect 18886 10013 18898 10016
rect 18840 10007 18898 10013
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 7616 9948 8064 9976
rect 7616 9936 7622 9948
rect 10594 9936 10600 9988
rect 10652 9976 10658 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 10652 9948 10701 9976
rect 10652 9936 10658 9948
rect 10689 9945 10701 9948
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 11146 9936 11152 9988
rect 11204 9936 11210 9988
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 12437 9979 12495 9985
rect 12437 9976 12449 9979
rect 12216 9948 12449 9976
rect 12216 9936 12222 9948
rect 12437 9945 12449 9948
rect 12483 9945 12495 9979
rect 12437 9939 12495 9945
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9945 15531 9979
rect 16022 9976 16028 9988
rect 15983 9948 16028 9976
rect 15473 9939 15531 9945
rect 10137 9911 10195 9917
rect 10137 9877 10149 9911
rect 10183 9908 10195 9911
rect 10318 9908 10324 9920
rect 10183 9880 10324 9908
rect 10183 9877 10195 9880
rect 10137 9871 10195 9877
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 15488 9908 15516 9939
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 16666 9976 16672 9988
rect 16627 9948 16672 9976
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 18690 9976 18696 9988
rect 16776 9948 18696 9976
rect 16776 9908 16804 9948
rect 18690 9936 18696 9948
rect 18748 9936 18754 9988
rect 22094 9976 22100 9988
rect 22055 9948 22100 9976
rect 22094 9936 22100 9948
rect 22152 9936 22158 9988
rect 15436 9880 16804 9908
rect 15436 9868 15442 9880
rect 19058 9868 19064 9920
rect 19116 9908 19122 9920
rect 19337 9911 19395 9917
rect 19337 9908 19349 9911
rect 19116 9880 19349 9908
rect 19116 9868 19122 9880
rect 19337 9877 19349 9880
rect 19383 9877 19395 9911
rect 19337 9871 19395 9877
rect 20070 9868 20076 9920
rect 20128 9908 20134 9920
rect 20257 9911 20315 9917
rect 20257 9908 20269 9911
rect 20128 9880 20269 9908
rect 20128 9868 20134 9880
rect 20257 9877 20269 9880
rect 20303 9877 20315 9911
rect 20257 9871 20315 9877
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22572 9908 22600 9976
rect 22060 9880 22600 9908
rect 22060 9868 22066 9880
rect 1104 9818 28336 9840
rect 1104 9766 1782 9818
rect 1834 9766 1846 9818
rect 1898 9766 1910 9818
rect 1962 9766 1974 9818
rect 2026 9766 4782 9818
rect 4834 9766 4846 9818
rect 4898 9766 4910 9818
rect 4962 9766 4974 9818
rect 5026 9766 7782 9818
rect 7834 9766 7846 9818
rect 7898 9766 7910 9818
rect 7962 9766 7974 9818
rect 8026 9766 10782 9818
rect 10834 9766 10846 9818
rect 10898 9766 10910 9818
rect 10962 9766 10974 9818
rect 11026 9766 13782 9818
rect 13834 9766 13846 9818
rect 13898 9766 13910 9818
rect 13962 9766 13974 9818
rect 14026 9766 16782 9818
rect 16834 9766 16846 9818
rect 16898 9766 16910 9818
rect 16962 9766 16974 9818
rect 17026 9766 19782 9818
rect 19834 9766 19846 9818
rect 19898 9766 19910 9818
rect 19962 9766 19974 9818
rect 20026 9766 22782 9818
rect 22834 9766 22846 9818
rect 22898 9766 22910 9818
rect 22962 9766 22974 9818
rect 23026 9766 25782 9818
rect 25834 9766 25846 9818
rect 25898 9766 25910 9818
rect 25962 9766 25974 9818
rect 26026 9766 28336 9818
rect 1104 9744 28336 9766
rect 5721 9707 5779 9713
rect 5721 9673 5733 9707
rect 5767 9704 5779 9707
rect 8294 9704 8300 9716
rect 5767 9676 8300 9704
rect 5767 9673 5779 9676
rect 5721 9667 5779 9673
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 8720 9676 9781 9704
rect 8720 9664 8726 9676
rect 9769 9673 9781 9676
rect 9815 9704 9827 9707
rect 10410 9704 10416 9716
rect 9815 9676 10416 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11204 9676 11805 9704
rect 11204 9664 11210 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 13630 9704 13636 9716
rect 11940 9676 13636 9704
rect 11940 9664 11946 9676
rect 13630 9664 13636 9676
rect 13688 9704 13694 9716
rect 14185 9707 14243 9713
rect 13688 9676 13814 9704
rect 13688 9664 13694 9676
rect 6089 9639 6147 9645
rect 6089 9605 6101 9639
rect 6135 9636 6147 9639
rect 6178 9636 6184 9648
rect 6135 9608 6184 9636
rect 6135 9605 6147 9608
rect 6089 9599 6147 9605
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 6457 9639 6515 9645
rect 6457 9605 6469 9639
rect 6503 9636 6515 9639
rect 7558 9636 7564 9648
rect 6503 9608 7564 9636
rect 6503 9605 6515 9608
rect 6457 9599 6515 9605
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 7742 9596 7748 9648
rect 7800 9596 7806 9648
rect 9401 9639 9459 9645
rect 9401 9605 9413 9639
rect 9447 9636 9459 9639
rect 9447 9608 10732 9636
rect 9447 9605 9459 9608
rect 9401 9599 9459 9605
rect 10502 9568 10508 9580
rect 10463 9540 10508 9568
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 10704 9577 10732 9608
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 13354 9636 13360 9648
rect 11296 9608 13360 9636
rect 11296 9596 11302 9608
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 13786 9636 13814 9676
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14918 9704 14924 9716
rect 14231 9676 14924 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 14918 9664 14924 9676
rect 14976 9664 14982 9716
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 21545 9707 21603 9713
rect 21545 9673 21557 9707
rect 21591 9704 21603 9707
rect 22002 9704 22008 9716
rect 21591 9676 22008 9704
rect 21591 9673 21603 9676
rect 21545 9667 21603 9673
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22094 9664 22100 9716
rect 22152 9704 22158 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 22152 9676 22661 9704
rect 22152 9664 22158 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 15013 9639 15071 9645
rect 15013 9636 15025 9639
rect 13786 9608 15025 9636
rect 15013 9605 15025 9608
rect 15059 9636 15071 9639
rect 16298 9636 16304 9648
rect 15059 9608 16304 9636
rect 15059 9605 15071 9608
rect 15013 9599 15071 9605
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 17494 9636 17500 9648
rect 16684 9608 17500 9636
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11514 9568 11520 9580
rect 11011 9540 11520 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 7006 9500 7012 9512
rect 6967 9472 7012 9500
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 7282 9500 7288 9512
rect 7243 9472 7288 9500
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9582 9500 9588 9512
rect 9079 9472 9588 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9500 10103 9503
rect 10594 9500 10600 9512
rect 10091 9472 10600 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10704 9500 10732 9531
rect 11514 9528 11520 9540
rect 11572 9568 11578 9580
rect 11882 9568 11888 9580
rect 11572 9540 11888 9568
rect 11572 9528 11578 9540
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 13127 9540 14381 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 14369 9537 14381 9540
rect 14415 9568 14427 9571
rect 14458 9568 14464 9580
rect 14415 9540 14464 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9568 15991 9571
rect 16114 9568 16120 9580
rect 15979 9540 16120 9568
rect 15979 9537 15991 9540
rect 15933 9531 15991 9537
rect 16114 9528 16120 9540
rect 16172 9568 16178 9580
rect 16485 9571 16543 9577
rect 16485 9568 16497 9571
rect 16172 9540 16497 9568
rect 16172 9528 16178 9540
rect 16485 9537 16497 9540
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16684 9577 16712 9608
rect 17494 9596 17500 9608
rect 17552 9636 17558 9648
rect 17681 9639 17739 9645
rect 17681 9636 17693 9639
rect 17552 9608 17693 9636
rect 17552 9596 17558 9608
rect 17681 9605 17693 9608
rect 17727 9636 17739 9639
rect 20257 9639 20315 9645
rect 17727 9608 19288 9636
rect 17727 9605 17739 9608
rect 17681 9599 17739 9605
rect 19260 9580 19288 9608
rect 20257 9605 20269 9639
rect 20303 9636 20315 9639
rect 21082 9636 21088 9648
rect 20303 9608 21088 9636
rect 20303 9605 20315 9608
rect 20257 9599 20315 9605
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16632 9540 16681 9568
rect 16632 9528 16638 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 19058 9568 19064 9580
rect 19019 9540 19064 9568
rect 18877 9531 18935 9537
rect 10778 9500 10784 9512
rect 10704 9472 10784 9500
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 11146 9500 11152 9512
rect 11107 9472 11152 9500
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9469 11483 9503
rect 11425 9463 11483 9469
rect 9122 9392 9128 9444
rect 9180 9432 9186 9444
rect 11440 9432 11468 9463
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 14182 9500 14188 9512
rect 13596 9472 14188 9500
rect 13596 9460 13602 9472
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 15838 9500 15844 9512
rect 15799 9472 15844 9500
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 18892 9500 18920 9531
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19242 9568 19248 9580
rect 19203 9540 19248 9568
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 19518 9528 19524 9580
rect 19576 9568 19582 9580
rect 20404 9571 20462 9577
rect 20404 9568 20416 9571
rect 19576 9540 20416 9568
rect 19576 9528 19582 9540
rect 20404 9537 20416 9540
rect 20450 9537 20462 9571
rect 21818 9568 21824 9580
rect 21779 9540 21824 9568
rect 20404 9531 20462 9537
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 23017 9571 23075 9577
rect 23017 9568 23029 9571
rect 21968 9540 23029 9568
rect 21968 9528 21974 9540
rect 23017 9537 23029 9540
rect 23063 9537 23075 9571
rect 23017 9531 23075 9537
rect 18966 9500 18972 9512
rect 18892 9472 18972 9500
rect 18966 9460 18972 9472
rect 19024 9460 19030 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 20088 9472 20637 9500
rect 9180 9404 11468 9432
rect 18693 9435 18751 9441
rect 9180 9392 9186 9404
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 19978 9432 19984 9444
rect 18739 9404 19984 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 19978 9392 19984 9404
rect 20036 9392 20042 9444
rect 20088 9376 20116 9472
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 22278 9500 22284 9512
rect 22239 9472 22284 9500
rect 20625 9463 20683 9469
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 20530 9432 20536 9444
rect 20491 9404 20536 9432
rect 20530 9392 20536 9404
rect 20588 9392 20594 9444
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 22186 9432 22192 9444
rect 21140 9404 22192 9432
rect 21140 9392 21146 9404
rect 22186 9392 22192 9404
rect 22244 9392 22250 9444
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 13412 9336 13461 9364
rect 13412 9324 13418 9336
rect 13449 9333 13461 9336
rect 13495 9364 13507 9367
rect 14182 9364 14188 9376
rect 13495 9336 14188 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 16945 9367 17003 9373
rect 16945 9333 16957 9367
rect 16991 9364 17003 9367
rect 17126 9364 17132 9376
rect 16991 9336 17132 9364
rect 16991 9333 17003 9336
rect 16945 9327 17003 9333
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 19797 9367 19855 9373
rect 19797 9333 19809 9367
rect 19843 9364 19855 9367
rect 20070 9364 20076 9376
rect 19843 9336 20076 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20901 9367 20959 9373
rect 20901 9333 20913 9367
rect 20947 9364 20959 9367
rect 21726 9364 21732 9376
rect 20947 9336 21732 9364
rect 20947 9333 20959 9336
rect 20901 9327 20959 9333
rect 21726 9324 21732 9336
rect 21784 9324 21790 9376
rect 1104 9274 28336 9296
rect 1104 9222 3282 9274
rect 3334 9222 3346 9274
rect 3398 9222 3410 9274
rect 3462 9222 3474 9274
rect 3526 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 6410 9274
rect 6462 9222 6474 9274
rect 6526 9222 9282 9274
rect 9334 9222 9346 9274
rect 9398 9222 9410 9274
rect 9462 9222 9474 9274
rect 9526 9222 12282 9274
rect 12334 9222 12346 9274
rect 12398 9222 12410 9274
rect 12462 9222 12474 9274
rect 12526 9222 15282 9274
rect 15334 9222 15346 9274
rect 15398 9222 15410 9274
rect 15462 9222 15474 9274
rect 15526 9222 18282 9274
rect 18334 9222 18346 9274
rect 18398 9222 18410 9274
rect 18462 9222 18474 9274
rect 18526 9222 21282 9274
rect 21334 9222 21346 9274
rect 21398 9222 21410 9274
rect 21462 9222 21474 9274
rect 21526 9222 24282 9274
rect 24334 9222 24346 9274
rect 24398 9222 24410 9274
rect 24462 9222 24474 9274
rect 24526 9222 27282 9274
rect 27334 9222 27346 9274
rect 27398 9222 27410 9274
rect 27462 9222 27474 9274
rect 27526 9222 28336 9274
rect 1104 9200 28336 9222
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 7653 9163 7711 9169
rect 7653 9160 7665 9163
rect 7340 9132 7665 9160
rect 7340 9120 7346 9132
rect 7653 9129 7665 9132
rect 7699 9129 7711 9163
rect 7653 9123 7711 9129
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8352 9132 8493 9160
rect 8352 9120 8358 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 8481 9123 8539 9129
rect 9122 9120 9128 9172
rect 9180 9160 9186 9172
rect 9217 9163 9275 9169
rect 9217 9160 9229 9163
rect 9180 9132 9229 9160
rect 9180 9120 9186 9132
rect 9217 9129 9229 9132
rect 9263 9129 9275 9163
rect 9217 9123 9275 9129
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10652 9132 10701 9160
rect 10652 9120 10658 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 10689 9123 10747 9129
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 11333 9163 11391 9169
rect 11333 9160 11345 9163
rect 10836 9132 11345 9160
rect 10836 9120 10842 9132
rect 11333 9129 11345 9132
rect 11379 9129 11391 9163
rect 11333 9123 11391 9129
rect 15841 9163 15899 9169
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 16114 9160 16120 9172
rect 15887 9132 16120 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 16574 9160 16580 9172
rect 16535 9132 16580 9160
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 19153 9163 19211 9169
rect 19153 9160 19165 9163
rect 18748 9132 19165 9160
rect 18748 9120 18754 9132
rect 19153 9129 19165 9132
rect 19199 9129 19211 9163
rect 19153 9123 19211 9129
rect 19242 9120 19248 9172
rect 19300 9160 19306 9172
rect 19889 9163 19947 9169
rect 19889 9160 19901 9163
rect 19300 9132 19901 9160
rect 19300 9120 19306 9132
rect 19889 9129 19901 9132
rect 19935 9129 19947 9163
rect 19889 9123 19947 9129
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22152 9132 22293 9160
rect 22152 9120 22158 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 6549 9095 6607 9101
rect 6549 9061 6561 9095
rect 6595 9092 6607 9095
rect 7009 9095 7067 9101
rect 7009 9092 7021 9095
rect 6595 9064 7021 9092
rect 6595 9061 6607 9064
rect 6549 9055 6607 9061
rect 7009 9061 7021 9064
rect 7055 9092 7067 9095
rect 7742 9092 7748 9104
rect 7055 9064 7748 9092
rect 7055 9061 7067 9064
rect 7009 9055 7067 9061
rect 7742 9052 7748 9064
rect 7800 9052 7806 9104
rect 21910 9052 21916 9104
rect 21968 9092 21974 9104
rect 22741 9095 22799 9101
rect 22741 9092 22753 9095
rect 21968 9064 22753 9092
rect 21968 9052 21974 9064
rect 22741 9061 22753 9064
rect 22787 9061 22799 9095
rect 22741 9055 22799 9061
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 7098 9024 7104 9036
rect 6788 8996 7104 9024
rect 6788 8984 6794 8996
rect 7098 8984 7104 8996
rect 7156 9024 7162 9036
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 7156 8996 7389 9024
rect 7156 8984 7162 8996
rect 7377 8993 7389 8996
rect 7423 9024 7435 9027
rect 8662 9024 8668 9036
rect 7423 8996 8668 9024
rect 7423 8993 7435 8996
rect 7377 8987 7435 8993
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 10502 9024 10508 9036
rect 10459 8996 10508 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 10502 8984 10508 8996
rect 10560 9024 10566 9036
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 10560 8996 11897 9024
rect 10560 8984 10566 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 9024 12771 9027
rect 13446 9024 13452 9036
rect 12759 8996 13452 9024
rect 12759 8993 12771 8996
rect 12713 8987 12771 8993
rect 13446 8984 13452 8996
rect 13504 9024 13510 9036
rect 13679 9027 13737 9033
rect 13679 9024 13691 9027
rect 13504 8996 13691 9024
rect 13504 8984 13510 8996
rect 13679 8993 13691 8996
rect 13725 8993 13737 9027
rect 13679 8987 13737 8993
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15838 9024 15844 9036
rect 14967 8996 15844 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 17126 9024 17132 9036
rect 17087 8996 17132 9024
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 18874 9024 18880 9036
rect 18835 8996 18880 9024
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 21082 9024 21088 9036
rect 21043 8996 21088 9024
rect 21082 8984 21088 8996
rect 21140 8984 21146 9036
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6144 8928 6837 8956
rect 6144 8916 6150 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8389 8959 8447 8965
rect 8389 8956 8401 8959
rect 8168 8928 8401 8956
rect 8168 8916 8174 8928
rect 8389 8925 8401 8928
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 8205 8891 8263 8897
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 9858 8888 9864 8900
rect 8251 8860 9864 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 10060 8888 10088 8919
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 10192 8928 11253 8956
rect 10192 8916 10198 8928
rect 11241 8925 11253 8928
rect 11287 8956 11299 8959
rect 12158 8956 12164 8968
rect 11287 8928 12164 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8956 13875 8959
rect 13863 8928 14412 8956
rect 13863 8925 13875 8928
rect 13817 8919 13875 8925
rect 10226 8888 10232 8900
rect 10060 8860 10232 8888
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 11057 8891 11115 8897
rect 11057 8857 11069 8891
rect 11103 8888 11115 8891
rect 11790 8888 11796 8900
rect 11103 8860 11796 8888
rect 11103 8857 11115 8860
rect 11057 8851 11115 8857
rect 11790 8848 11796 8860
rect 11848 8848 11854 8900
rect 12989 8891 13047 8897
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13170 8888 13176 8900
rect 13035 8860 13176 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13170 8848 13176 8860
rect 13228 8848 13234 8900
rect 6178 8820 6184 8832
rect 6139 8792 6184 8820
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 14384 8829 14412 8928
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16724 8928 16865 8956
rect 16724 8916 16730 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 19150 8916 19156 8968
rect 19208 8956 19214 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19208 8928 19717 8956
rect 19208 8916 19214 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 21266 8956 21272 8968
rect 20036 8928 21272 8956
rect 20036 8916 20042 8928
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 21692 8928 21741 8956
rect 21692 8916 21698 8928
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8956 21879 8959
rect 22278 8956 22284 8968
rect 21867 8928 22284 8956
rect 21867 8925 21879 8928
rect 21821 8919 21879 8925
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 17678 8848 17684 8900
rect 17736 8848 17742 8900
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 20714 8888 20720 8900
rect 19392 8860 20720 8888
rect 19392 8848 19398 8860
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 22186 8848 22192 8900
rect 22244 8888 22250 8900
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 22244 8860 23121 8888
rect 22244 8848 22250 8860
rect 23109 8857 23121 8860
rect 23155 8857 23167 8891
rect 23109 8851 23167 8857
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8820 14427 8823
rect 14458 8820 14464 8832
rect 14415 8792 14464 8820
rect 14415 8789 14427 8792
rect 14369 8783 14427 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20257 8823 20315 8829
rect 20257 8820 20269 8823
rect 20128 8792 20269 8820
rect 20128 8780 20134 8792
rect 20257 8789 20269 8792
rect 20303 8789 20315 8823
rect 20257 8783 20315 8789
rect 1104 8730 28336 8752
rect 1104 8678 1782 8730
rect 1834 8678 1846 8730
rect 1898 8678 1910 8730
rect 1962 8678 1974 8730
rect 2026 8678 4782 8730
rect 4834 8678 4846 8730
rect 4898 8678 4910 8730
rect 4962 8678 4974 8730
rect 5026 8678 7782 8730
rect 7834 8678 7846 8730
rect 7898 8678 7910 8730
rect 7962 8678 7974 8730
rect 8026 8678 10782 8730
rect 10834 8678 10846 8730
rect 10898 8678 10910 8730
rect 10962 8678 10974 8730
rect 11026 8678 13782 8730
rect 13834 8678 13846 8730
rect 13898 8678 13910 8730
rect 13962 8678 13974 8730
rect 14026 8678 16782 8730
rect 16834 8678 16846 8730
rect 16898 8678 16910 8730
rect 16962 8678 16974 8730
rect 17026 8678 19782 8730
rect 19834 8678 19846 8730
rect 19898 8678 19910 8730
rect 19962 8678 19974 8730
rect 20026 8678 22782 8730
rect 22834 8678 22846 8730
rect 22898 8678 22910 8730
rect 22962 8678 22974 8730
rect 23026 8678 25782 8730
rect 25834 8678 25846 8730
rect 25898 8678 25910 8730
rect 25962 8678 25974 8730
rect 26026 8678 28336 8730
rect 1104 8656 28336 8678
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 7374 8616 7380 8628
rect 6135 8588 7380 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 7374 8576 7380 8588
rect 7432 8616 7438 8628
rect 8110 8616 8116 8628
rect 7432 8588 8116 8616
rect 7432 8576 7438 8588
rect 8110 8576 8116 8588
rect 8168 8616 8174 8628
rect 8754 8616 8760 8628
rect 8168 8588 8760 8616
rect 8168 8576 8174 8588
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 11514 8616 11520 8628
rect 10551 8588 11520 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 16666 8616 16672 8628
rect 13412 8588 16672 8616
rect 13412 8576 13418 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 17184 8588 17233 8616
rect 17184 8576 17190 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17678 8616 17684 8628
rect 17639 8588 17684 8616
rect 17221 8579 17279 8585
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 18417 8619 18475 8625
rect 18417 8585 18429 8619
rect 18463 8616 18475 8619
rect 18598 8616 18604 8628
rect 18463 8588 18604 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 18598 8576 18604 8588
rect 18656 8616 18662 8628
rect 18782 8616 18788 8628
rect 18656 8588 18788 8616
rect 18656 8576 18662 8588
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 19061 8619 19119 8625
rect 19061 8585 19073 8619
rect 19107 8616 19119 8619
rect 19150 8616 19156 8628
rect 19107 8588 19156 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 20530 8576 20536 8628
rect 20588 8616 20594 8628
rect 21174 8616 21180 8628
rect 20588 8588 21180 8616
rect 20588 8576 20594 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 21266 8576 21272 8628
rect 21324 8616 21330 8628
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 21324 8588 21557 8616
rect 21324 8576 21330 8588
rect 21545 8585 21557 8588
rect 21591 8616 21603 8619
rect 21818 8616 21824 8628
rect 21591 8588 21824 8616
rect 21591 8585 21603 8588
rect 21545 8579 21603 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 22649 8619 22707 8625
rect 22649 8616 22661 8619
rect 22244 8588 22661 8616
rect 22244 8576 22250 8588
rect 22649 8585 22661 8588
rect 22695 8585 22707 8619
rect 22649 8579 22707 8585
rect 7650 8548 7656 8560
rect 7611 8520 7656 8548
rect 7650 8508 7656 8520
rect 7708 8508 7714 8560
rect 8021 8551 8079 8557
rect 8021 8517 8033 8551
rect 8067 8548 8079 8551
rect 8481 8551 8539 8557
rect 8481 8548 8493 8551
rect 8067 8520 8493 8548
rect 8067 8517 8079 8520
rect 8021 8511 8079 8517
rect 8481 8517 8493 8520
rect 8527 8548 8539 8551
rect 8570 8548 8576 8560
rect 8527 8520 8576 8548
rect 8527 8517 8539 8520
rect 8481 8511 8539 8517
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 10042 8548 10048 8560
rect 9324 8520 10048 8548
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8480 7251 8483
rect 8294 8480 8300 8492
rect 7239 8452 8300 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 9324 8489 9352 8520
rect 10042 8508 10048 8520
rect 10100 8548 10106 8560
rect 11808 8548 11836 8576
rect 10100 8520 11836 8548
rect 10100 8508 10106 8520
rect 13630 8508 13636 8560
rect 13688 8508 13694 8560
rect 14458 8508 14464 8560
rect 14516 8548 14522 8560
rect 14921 8551 14979 8557
rect 14921 8548 14933 8551
rect 14516 8520 14933 8548
rect 14516 8508 14522 8520
rect 14921 8517 14933 8520
rect 14967 8517 14979 8551
rect 14921 8511 14979 8517
rect 15381 8551 15439 8557
rect 15381 8517 15393 8551
rect 15427 8548 15439 8551
rect 15654 8548 15660 8560
rect 15427 8520 15660 8548
rect 15427 8517 15439 8520
rect 15381 8511 15439 8517
rect 15654 8508 15660 8520
rect 15712 8548 15718 8560
rect 19168 8548 19196 8576
rect 20438 8548 20444 8560
rect 15712 8520 17816 8548
rect 19168 8520 20444 8548
rect 15712 8508 15718 8520
rect 17788 8492 17816 8520
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 11422 8480 11428 8492
rect 9309 8443 9367 8449
rect 9416 8452 11100 8480
rect 11383 8452 11428 8480
rect 7098 8412 7104 8424
rect 7059 8384 7104 8412
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 9030 8412 9036 8424
rect 8943 8384 9036 8412
rect 9030 8372 9036 8384
rect 9088 8412 9094 8424
rect 9416 8412 9444 8452
rect 9088 8384 9444 8412
rect 9493 8415 9551 8421
rect 9088 8372 9094 8384
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9582 8412 9588 8424
rect 9539 8384 9588 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 10778 8412 10784 8424
rect 10739 8384 10784 8412
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 11072 8412 11100 8452
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 15838 8480 15844 8492
rect 15799 8452 15844 8480
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 17770 8440 17776 8492
rect 17828 8480 17834 8492
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 17828 8452 18245 8480
rect 17828 8440 17834 8452
rect 18233 8449 18245 8452
rect 18279 8480 18291 8483
rect 18874 8480 18880 8492
rect 18279 8452 18880 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 11238 8412 11244 8424
rect 11072 8384 11244 8412
rect 11238 8372 11244 8384
rect 11296 8412 11302 8424
rect 11974 8412 11980 8424
rect 11296 8384 11980 8412
rect 11296 8372 11302 8384
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12894 8412 12900 8424
rect 12855 8384 12900 8412
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 13170 8412 13176 8424
rect 13131 8384 13176 8412
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 7616 8316 10057 8344
rect 7616 8304 7622 8316
rect 10045 8313 10057 8316
rect 10091 8344 10103 8347
rect 11146 8344 11152 8356
rect 10091 8316 11152 8344
rect 10091 8313 10103 8316
rect 10045 8307 10103 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 16945 8347 17003 8353
rect 16945 8344 16957 8347
rect 16724 8316 16957 8344
rect 16724 8304 16730 8316
rect 16945 8313 16957 8316
rect 16991 8344 17003 8347
rect 19334 8344 19340 8356
rect 16991 8316 19340 8344
rect 16991 8313 17003 8316
rect 16945 8307 17003 8313
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 19444 8344 19472 8443
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19702 8480 19708 8492
rect 19576 8452 19621 8480
rect 19663 8452 19708 8480
rect 19576 8440 19582 8452
rect 19702 8440 19708 8452
rect 19760 8440 19766 8492
rect 20088 8489 20116 8520
rect 20438 8508 20444 8520
rect 20496 8548 20502 8560
rect 22002 8548 22008 8560
rect 20496 8520 22008 8548
rect 20496 8508 20502 8520
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8449 20131 8483
rect 20266 8483 20324 8489
rect 20266 8480 20278 8483
rect 20073 8443 20131 8449
rect 20180 8452 20278 8480
rect 20070 8344 20076 8356
rect 19444 8316 20076 8344
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 20180 8344 20208 8452
rect 20266 8449 20278 8452
rect 20312 8449 20324 8483
rect 20266 8443 20324 8449
rect 21634 8440 21640 8492
rect 21692 8480 21698 8492
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 21692 8452 21925 8480
rect 21692 8440 21698 8452
rect 21913 8449 21925 8452
rect 21959 8449 21971 8483
rect 21913 8443 21971 8449
rect 20622 8412 20628 8424
rect 20583 8384 20628 8412
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 22462 8344 22468 8356
rect 20180 8316 22468 8344
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 6144 8248 6377 8276
rect 6144 8236 6150 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 11164 8276 11192 8304
rect 14550 8276 14556 8288
rect 11164 8248 14556 8276
rect 6365 8239 6423 8245
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 16209 8279 16267 8285
rect 16209 8245 16221 8279
rect 16255 8276 16267 8279
rect 16298 8276 16304 8288
rect 16255 8248 16304 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 19242 8236 19248 8288
rect 19300 8276 19306 8288
rect 20180 8276 20208 8316
rect 22462 8304 22468 8316
rect 22520 8304 22526 8356
rect 22278 8276 22284 8288
rect 19300 8248 20208 8276
rect 22239 8248 22284 8276
rect 19300 8236 19306 8248
rect 22278 8236 22284 8248
rect 22336 8236 22342 8288
rect 1104 8186 28336 8208
rect 1104 8134 3282 8186
rect 3334 8134 3346 8186
rect 3398 8134 3410 8186
rect 3462 8134 3474 8186
rect 3526 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 6410 8186
rect 6462 8134 6474 8186
rect 6526 8134 9282 8186
rect 9334 8134 9346 8186
rect 9398 8134 9410 8186
rect 9462 8134 9474 8186
rect 9526 8134 12282 8186
rect 12334 8134 12346 8186
rect 12398 8134 12410 8186
rect 12462 8134 12474 8186
rect 12526 8134 15282 8186
rect 15334 8134 15346 8186
rect 15398 8134 15410 8186
rect 15462 8134 15474 8186
rect 15526 8134 18282 8186
rect 18334 8134 18346 8186
rect 18398 8134 18410 8186
rect 18462 8134 18474 8186
rect 18526 8134 21282 8186
rect 21334 8134 21346 8186
rect 21398 8134 21410 8186
rect 21462 8134 21474 8186
rect 21526 8134 24282 8186
rect 24334 8134 24346 8186
rect 24398 8134 24410 8186
rect 24462 8134 24474 8186
rect 24526 8134 27282 8186
rect 27334 8134 27346 8186
rect 27398 8134 27410 8186
rect 27462 8134 27474 8186
rect 27526 8134 28336 8186
rect 1104 8112 28336 8134
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 9030 8072 9036 8084
rect 8991 8044 9036 8072
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 10226 8072 10232 8084
rect 9180 8044 10232 8072
rect 9180 8032 9186 8044
rect 10226 8032 10232 8044
rect 10284 8072 10290 8084
rect 11241 8075 11299 8081
rect 11241 8072 11253 8075
rect 10284 8044 11253 8072
rect 10284 8032 10290 8044
rect 11241 8041 11253 8044
rect 11287 8041 11299 8075
rect 11241 8035 11299 8041
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13170 8072 13176 8084
rect 13035 8044 13176 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13504 8044 14197 8072
rect 13504 8032 13510 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 14185 8035 14243 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16206 8072 16212 8084
rect 16167 8044 16212 8072
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 17865 8075 17923 8081
rect 17865 8041 17877 8075
rect 17911 8072 17923 8075
rect 19058 8072 19064 8084
rect 17911 8044 19064 8072
rect 17911 8041 17923 8044
rect 17865 8035 17923 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 22278 8072 22284 8084
rect 21407 8044 22284 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 10134 8004 10140 8016
rect 8812 7976 10140 8004
rect 8812 7964 8818 7976
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10965 8007 11023 8013
rect 10965 7973 10977 8007
rect 11011 8004 11023 8007
rect 11422 8004 11428 8016
rect 11011 7976 11428 8004
rect 11011 7973 11023 7976
rect 10965 7967 11023 7973
rect 11422 7964 11428 7976
rect 11480 8004 11486 8016
rect 18325 8007 18383 8013
rect 18325 8004 18337 8007
rect 11480 7976 18337 8004
rect 11480 7964 11486 7976
rect 18325 7973 18337 7976
rect 18371 8004 18383 8007
rect 19702 8004 19708 8016
rect 18371 7976 19708 8004
rect 18371 7973 18383 7976
rect 18325 7967 18383 7973
rect 19702 7964 19708 7976
rect 19760 8004 19766 8016
rect 20806 8004 20812 8016
rect 19760 7976 20812 8004
rect 19760 7964 19766 7976
rect 20806 7964 20812 7976
rect 20864 8004 20870 8016
rect 20864 7976 21588 8004
rect 20864 7964 20870 7976
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7936 6883 7939
rect 8294 7936 8300 7948
rect 6871 7908 8300 7936
rect 6871 7905 6883 7908
rect 6825 7899 6883 7905
rect 8294 7896 8300 7908
rect 8352 7936 8358 7948
rect 10778 7936 10784 7948
rect 8352 7908 10784 7936
rect 8352 7896 8358 7908
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 13817 7939 13875 7945
rect 13817 7936 13829 7939
rect 13596 7908 13829 7936
rect 13596 7896 13602 7908
rect 13817 7905 13829 7908
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 16022 7896 16028 7948
rect 16080 7936 16086 7948
rect 18693 7939 18751 7945
rect 16080 7908 18184 7936
rect 16080 7896 16086 7908
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6236 7840 6469 7868
rect 6236 7828 6242 7840
rect 6457 7837 6469 7840
rect 6503 7868 6515 7871
rect 7006 7868 7012 7880
rect 6503 7840 7012 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 7006 7828 7012 7840
rect 7064 7868 7070 7880
rect 8573 7871 8631 7877
rect 8573 7868 8585 7871
rect 7064 7840 8585 7868
rect 7064 7828 7070 7840
rect 8573 7837 8585 7840
rect 8619 7837 8631 7871
rect 8754 7868 8760 7880
rect 8715 7840 8760 7868
rect 8573 7831 8631 7837
rect 7466 7760 7472 7812
rect 7524 7800 7530 7812
rect 7745 7803 7803 7809
rect 7745 7800 7757 7803
rect 7524 7772 7757 7800
rect 7524 7760 7530 7772
rect 7745 7769 7757 7772
rect 7791 7769 7803 7803
rect 8588 7800 8616 7831
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 9640 7840 9873 7868
rect 9640 7828 9646 7840
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 9600 7800 9628 7828
rect 8588 7772 9628 7800
rect 9876 7800 9904 7831
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10134 7868 10140 7880
rect 10008 7840 10053 7868
rect 10095 7840 10140 7868
rect 10008 7828 10014 7840
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 10376 7840 12541 7868
rect 10376 7828 10382 7840
rect 12529 7837 12541 7840
rect 12575 7868 12587 7871
rect 13354 7868 13360 7880
rect 12575 7840 12848 7868
rect 13315 7840 13360 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 10226 7800 10232 7812
rect 9876 7772 10232 7800
rect 7745 7763 7803 7769
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 10597 7803 10655 7809
rect 10597 7769 10609 7803
rect 10643 7800 10655 7803
rect 12710 7800 12716 7812
rect 10643 7772 12716 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11572 7704 11621 7732
rect 11572 7692 11578 7704
rect 11609 7701 11621 7704
rect 11655 7701 11667 7735
rect 12250 7732 12256 7744
rect 12211 7704 12256 7732
rect 11609 7695 11667 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12820 7732 12848 7840
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 16666 7868 16672 7880
rect 16627 7840 16672 7868
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 18156 7877 18184 7908
rect 18693 7905 18705 7939
rect 18739 7936 18751 7939
rect 19150 7936 19156 7948
rect 18739 7908 19156 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 21560 7945 21588 7976
rect 21545 7939 21603 7945
rect 21545 7905 21557 7939
rect 21591 7905 21603 7939
rect 22002 7936 22008 7948
rect 21963 7908 22008 7936
rect 21545 7899 21603 7905
rect 22002 7896 22008 7908
rect 22060 7896 22066 7948
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18230 7868 18236 7880
rect 18187 7840 18236 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 18969 7871 19027 7877
rect 18969 7868 18981 7871
rect 18555 7840 18981 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 18969 7837 18981 7840
rect 19015 7868 19027 7871
rect 19518 7868 19524 7880
rect 19015 7840 19524 7868
rect 19015 7837 19027 7840
rect 18969 7831 19027 7837
rect 19518 7828 19524 7840
rect 19576 7868 19582 7880
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 19576 7840 20453 7868
rect 19576 7828 19582 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 21726 7868 21732 7880
rect 21687 7840 21732 7868
rect 20441 7831 20499 7837
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 17313 7803 17371 7809
rect 17313 7769 17325 7803
rect 17359 7800 17371 7803
rect 18690 7800 18696 7812
rect 17359 7772 18696 7800
rect 17359 7769 17371 7772
rect 17313 7763 17371 7769
rect 18690 7760 18696 7772
rect 18748 7760 18754 7812
rect 21174 7760 21180 7812
rect 21232 7800 21238 7812
rect 22112 7800 22140 7831
rect 21232 7772 22140 7800
rect 21232 7760 21238 7772
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 12820 7704 13553 7732
rect 13541 7701 13553 7704
rect 13587 7732 13599 7735
rect 13630 7732 13636 7744
rect 13587 7704 13636 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 16298 7692 16304 7744
rect 16356 7732 16362 7744
rect 18509 7735 18567 7741
rect 18509 7732 18521 7735
rect 16356 7704 18521 7732
rect 16356 7692 16362 7704
rect 18509 7701 18521 7704
rect 18555 7701 18567 7735
rect 18509 7695 18567 7701
rect 19242 7692 19248 7744
rect 19300 7732 19306 7744
rect 19337 7735 19395 7741
rect 19337 7732 19349 7735
rect 19300 7704 19349 7732
rect 19300 7692 19306 7704
rect 19337 7701 19349 7704
rect 19383 7701 19395 7735
rect 20070 7732 20076 7744
rect 20031 7704 20076 7732
rect 19337 7695 19395 7701
rect 20070 7692 20076 7704
rect 20128 7692 20134 7744
rect 1104 7642 28336 7664
rect 1104 7590 1782 7642
rect 1834 7590 1846 7642
rect 1898 7590 1910 7642
rect 1962 7590 1974 7642
rect 2026 7590 4782 7642
rect 4834 7590 4846 7642
rect 4898 7590 4910 7642
rect 4962 7590 4974 7642
rect 5026 7590 7782 7642
rect 7834 7590 7846 7642
rect 7898 7590 7910 7642
rect 7962 7590 7974 7642
rect 8026 7590 10782 7642
rect 10834 7590 10846 7642
rect 10898 7590 10910 7642
rect 10962 7590 10974 7642
rect 11026 7590 13782 7642
rect 13834 7590 13846 7642
rect 13898 7590 13910 7642
rect 13962 7590 13974 7642
rect 14026 7590 16782 7642
rect 16834 7590 16846 7642
rect 16898 7590 16910 7642
rect 16962 7590 16974 7642
rect 17026 7590 19782 7642
rect 19834 7590 19846 7642
rect 19898 7590 19910 7642
rect 19962 7590 19974 7642
rect 20026 7590 22782 7642
rect 22834 7590 22846 7642
rect 22898 7590 22910 7642
rect 22962 7590 22974 7642
rect 23026 7590 25782 7642
rect 25834 7590 25846 7642
rect 25898 7590 25910 7642
rect 25962 7590 25974 7642
rect 26026 7590 28336 7642
rect 1104 7568 28336 7590
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7374 7528 7380 7540
rect 7335 7500 7380 7528
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 7837 7531 7895 7537
rect 7837 7497 7849 7531
rect 7883 7528 7895 7531
rect 8294 7528 8300 7540
rect 7883 7500 8300 7528
rect 7883 7497 7895 7500
rect 7837 7491 7895 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 9916 7500 10057 7528
rect 9916 7488 9922 7500
rect 10045 7497 10057 7500
rect 10091 7497 10103 7531
rect 10045 7491 10103 7497
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 10284 7500 11621 7528
rect 10284 7488 10290 7500
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11609 7491 11667 7497
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13412 7500 13553 7528
rect 13412 7488 13418 7500
rect 13541 7497 13553 7500
rect 13587 7528 13599 7531
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13587 7500 13645 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 16666 7528 16672 7540
rect 16627 7500 16672 7528
rect 13633 7491 13691 7497
rect 16666 7488 16672 7500
rect 16724 7488 16730 7540
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 17359 7500 17693 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 17681 7497 17693 7500
rect 17727 7528 17739 7531
rect 17770 7528 17776 7540
rect 17727 7500 17776 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18230 7528 18236 7540
rect 18191 7500 18236 7528
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 20438 7528 20444 7540
rect 20399 7500 20444 7528
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 21726 7488 21732 7540
rect 21784 7528 21790 7540
rect 22189 7531 22247 7537
rect 22189 7528 22201 7531
rect 21784 7500 22201 7528
rect 21784 7488 21790 7500
rect 22189 7497 22201 7500
rect 22235 7497 22247 7531
rect 22189 7491 22247 7497
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 8481 7463 8539 7469
rect 8481 7460 8493 7463
rect 7156 7432 8493 7460
rect 7156 7420 7162 7432
rect 8481 7429 8493 7432
rect 8527 7460 8539 7463
rect 9677 7463 9735 7469
rect 9677 7460 9689 7463
rect 8527 7432 9689 7460
rect 8527 7429 8539 7432
rect 8481 7423 8539 7429
rect 9677 7429 9689 7432
rect 9723 7460 9735 7463
rect 9950 7460 9956 7472
rect 9723 7432 9956 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 10134 7420 10140 7472
rect 10192 7460 10198 7472
rect 11241 7463 11299 7469
rect 11241 7460 11253 7463
rect 10192 7432 11253 7460
rect 10192 7420 10198 7432
rect 11241 7429 11253 7432
rect 11287 7460 11299 7463
rect 11514 7460 11520 7472
rect 11287 7432 11520 7460
rect 11287 7429 11299 7432
rect 11241 7423 11299 7429
rect 11514 7420 11520 7432
rect 11572 7420 11578 7472
rect 12250 7420 12256 7472
rect 12308 7460 12314 7472
rect 12621 7463 12679 7469
rect 12621 7460 12633 7463
rect 12308 7432 12633 7460
rect 12308 7420 12314 7432
rect 12621 7429 12633 7432
rect 12667 7460 12679 7463
rect 12894 7460 12900 7472
rect 12667 7432 12900 7460
rect 12667 7429 12679 7432
rect 12621 7423 12679 7429
rect 12894 7420 12900 7432
rect 12952 7420 12958 7472
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 21174 7460 21180 7472
rect 14608 7432 15240 7460
rect 21135 7432 21180 7460
rect 14608 7420 14614 7432
rect 9122 7392 9128 7404
rect 9083 7364 9128 7392
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7361 10471 7395
rect 13262 7392 13268 7404
rect 13223 7364 13268 7392
rect 10413 7355 10471 7361
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 10318 7324 10324 7336
rect 6144 7296 10324 7324
rect 6144 7284 6150 7296
rect 10318 7284 10324 7296
rect 10376 7324 10382 7336
rect 10428 7324 10456 7355
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 14734 7392 14740 7404
rect 13596 7364 13814 7392
rect 14695 7364 14740 7392
rect 13596 7352 13602 7364
rect 10870 7324 10876 7336
rect 10376 7296 10876 7324
rect 10376 7284 10382 7296
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 13786 7324 13814 7364
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 15212 7401 15240 7432
rect 21174 7420 21180 7432
rect 21232 7420 21238 7472
rect 15197 7395 15255 7401
rect 14884 7364 14929 7392
rect 14884 7352 14890 7364
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 16114 7392 16120 7404
rect 15344 7364 16120 7392
rect 15344 7352 15350 7364
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7392 19119 7395
rect 19426 7392 19432 7404
rect 19107 7364 19432 7392
rect 19107 7361 19119 7364
rect 19061 7355 19119 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 22002 7392 22008 7404
rect 21867 7364 22008 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 22002 7352 22008 7364
rect 22060 7352 22066 7404
rect 14844 7324 14872 7352
rect 19334 7324 19340 7336
rect 13786 7296 14872 7324
rect 19295 7296 19340 7324
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 21726 7324 21732 7336
rect 19935 7296 21732 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 21726 7284 21732 7296
rect 21784 7284 21790 7336
rect 14274 7256 14280 7268
rect 13786 7228 14280 7256
rect 8205 7191 8263 7197
rect 8205 7157 8217 7191
rect 8251 7188 8263 7191
rect 10042 7188 10048 7200
rect 8251 7160 10048 7188
rect 8251 7157 8263 7160
rect 8205 7151 8263 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10594 7188 10600 7200
rect 10555 7160 10600 7188
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11146 7188 11152 7200
rect 11011 7160 11152 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 12066 7188 12072 7200
rect 12027 7160 12072 7188
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 13541 7191 13599 7197
rect 13541 7157 13553 7191
rect 13587 7188 13599 7191
rect 13786 7188 13814 7228
rect 14274 7216 14280 7228
rect 14332 7216 14338 7268
rect 14918 7216 14924 7268
rect 14976 7256 14982 7268
rect 19242 7256 19248 7268
rect 14976 7228 19248 7256
rect 14976 7216 14982 7228
rect 19242 7216 19248 7228
rect 19300 7216 19306 7268
rect 13587 7160 13814 7188
rect 14185 7191 14243 7197
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 14185 7157 14197 7191
rect 14231 7188 14243 7191
rect 14366 7188 14372 7200
rect 14231 7160 14372 7188
rect 14231 7157 14243 7160
rect 14185 7151 14243 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 16114 7188 16120 7200
rect 15795 7160 16120 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 18693 7191 18751 7197
rect 18693 7157 18705 7191
rect 18739 7188 18751 7191
rect 18966 7188 18972 7200
rect 18739 7160 18972 7188
rect 18739 7157 18751 7160
rect 18693 7151 18751 7157
rect 18966 7148 18972 7160
rect 19024 7188 19030 7200
rect 19610 7188 19616 7200
rect 19024 7160 19616 7188
rect 19024 7148 19030 7160
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 1104 7098 28336 7120
rect 1104 7046 3282 7098
rect 3334 7046 3346 7098
rect 3398 7046 3410 7098
rect 3462 7046 3474 7098
rect 3526 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 6410 7098
rect 6462 7046 6474 7098
rect 6526 7046 9282 7098
rect 9334 7046 9346 7098
rect 9398 7046 9410 7098
rect 9462 7046 9474 7098
rect 9526 7046 12282 7098
rect 12334 7046 12346 7098
rect 12398 7046 12410 7098
rect 12462 7046 12474 7098
rect 12526 7046 15282 7098
rect 15334 7046 15346 7098
rect 15398 7046 15410 7098
rect 15462 7046 15474 7098
rect 15526 7046 18282 7098
rect 18334 7046 18346 7098
rect 18398 7046 18410 7098
rect 18462 7046 18474 7098
rect 18526 7046 21282 7098
rect 21334 7046 21346 7098
rect 21398 7046 21410 7098
rect 21462 7046 21474 7098
rect 21526 7046 24282 7098
rect 24334 7046 24346 7098
rect 24398 7046 24410 7098
rect 24462 7046 24474 7098
rect 24526 7046 27282 7098
rect 27334 7046 27346 7098
rect 27398 7046 27410 7098
rect 27462 7046 27474 7098
rect 27526 7046 28336 7098
rect 1104 7024 28336 7046
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 9309 6987 9367 6993
rect 9309 6984 9321 6987
rect 8435 6956 9321 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 9309 6953 9321 6956
rect 9355 6984 9367 6987
rect 9858 6984 9864 6996
rect 9355 6956 9864 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 9858 6944 9864 6956
rect 9916 6984 9922 6996
rect 10137 6987 10195 6993
rect 10137 6984 10149 6987
rect 9916 6956 10149 6984
rect 9916 6944 9922 6956
rect 10137 6953 10149 6956
rect 10183 6953 10195 6987
rect 10870 6984 10876 6996
rect 10831 6956 10876 6984
rect 10137 6947 10195 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11790 6984 11796 6996
rect 11440 6956 11796 6984
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 9122 6916 9128 6928
rect 8803 6888 9128 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 7466 6780 7472 6792
rect 7427 6752 7472 6780
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7650 6780 7656 6792
rect 7611 6752 7656 6780
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8772 6780 8800 6879
rect 9122 6876 9128 6888
rect 9180 6876 9186 6928
rect 11440 6857 11468 6956
rect 11790 6944 11796 6956
rect 11848 6984 11854 6996
rect 13262 6984 13268 6996
rect 11848 6956 13268 6984
rect 11848 6944 11854 6956
rect 13262 6944 13268 6956
rect 13320 6984 13326 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13320 6956 13737 6984
rect 13320 6944 13326 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 14550 6984 14556 6996
rect 14511 6956 14556 6984
rect 13725 6947 13783 6953
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 14734 6944 14740 6996
rect 14792 6984 14798 6996
rect 16298 6984 16304 6996
rect 14792 6956 16304 6984
rect 14792 6944 14798 6956
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 16666 6944 16672 6996
rect 16724 6984 16730 6996
rect 16853 6987 16911 6993
rect 16853 6984 16865 6987
rect 16724 6956 16865 6984
rect 16724 6944 16730 6956
rect 16853 6953 16865 6956
rect 16899 6953 16911 6987
rect 16853 6947 16911 6953
rect 17678 6944 17684 6996
rect 17736 6984 17742 6996
rect 17865 6987 17923 6993
rect 17865 6984 17877 6987
rect 17736 6956 17877 6984
rect 17736 6944 17742 6956
rect 17865 6953 17877 6956
rect 17911 6953 17923 6987
rect 21174 6984 21180 6996
rect 21135 6956 21180 6984
rect 17865 6947 17923 6953
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 14277 6919 14335 6925
rect 14277 6885 14289 6919
rect 14323 6916 14335 6919
rect 15102 6916 15108 6928
rect 14323 6888 15108 6916
rect 14323 6885 14335 6888
rect 14277 6879 14335 6885
rect 15102 6876 15108 6888
rect 15160 6876 15166 6928
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6817 11483 6851
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 11425 6811 11483 6817
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15473 6851 15531 6857
rect 15473 6848 15485 6851
rect 14884 6820 15485 6848
rect 14884 6808 14890 6820
rect 15473 6817 15485 6820
rect 15519 6848 15531 6851
rect 15654 6848 15660 6860
rect 15519 6820 15660 6848
rect 15519 6817 15531 6820
rect 15473 6811 15531 6817
rect 15654 6808 15660 6820
rect 15712 6848 15718 6860
rect 16684 6848 16712 6944
rect 15712 6820 16712 6848
rect 19981 6851 20039 6857
rect 15712 6808 15718 6820
rect 19981 6817 19993 6851
rect 20027 6848 20039 6851
rect 20070 6848 20076 6860
rect 20027 6820 20076 6848
rect 20027 6817 20039 6820
rect 19981 6811 20039 6817
rect 20070 6808 20076 6820
rect 20128 6808 20134 6860
rect 10042 6780 10048 6792
rect 8067 6752 8800 6780
rect 10003 6752 10048 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 6822 6672 6828 6724
rect 6880 6712 6886 6724
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6880 6684 7021 6712
rect 6880 6672 6886 6684
rect 7009 6681 7021 6684
rect 7055 6712 7067 6715
rect 8036 6712 8064 6743
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 15565 6783 15623 6789
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 15838 6780 15844 6792
rect 15611 6752 15844 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 16666 6780 16672 6792
rect 16627 6752 16672 6780
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6780 17739 6783
rect 18138 6780 18144 6792
rect 17727 6752 18144 6780
rect 17727 6749 17739 6752
rect 17681 6743 17739 6749
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18601 6783 18659 6789
rect 18601 6749 18613 6783
rect 18647 6780 18659 6783
rect 19426 6780 19432 6792
rect 18647 6752 19432 6780
rect 18647 6749 18659 6752
rect 18601 6743 18659 6749
rect 19426 6740 19432 6752
rect 19484 6780 19490 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19484 6752 19901 6780
rect 19484 6740 19490 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 11698 6712 11704 6724
rect 7055 6684 8064 6712
rect 11659 6684 11704 6712
rect 7055 6681 7067 6684
rect 7009 6675 7067 6681
rect 11698 6672 11704 6684
rect 11756 6672 11762 6724
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 15930 6672 15936 6724
rect 15988 6712 15994 6724
rect 16025 6715 16083 6721
rect 16025 6712 16037 6715
rect 15988 6684 16037 6712
rect 15988 6672 15994 6684
rect 16025 6681 16037 6684
rect 16071 6681 16083 6715
rect 16025 6675 16083 6681
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6638 6644 6644 6656
rect 6503 6616 6644 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18877 6647 18935 6653
rect 18877 6644 18889 6647
rect 18012 6616 18889 6644
rect 18012 6604 18018 6616
rect 18877 6613 18889 6616
rect 18923 6644 18935 6647
rect 19334 6644 19340 6656
rect 18923 6616 19340 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19904 6644 19932 6743
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 21453 6783 21511 6789
rect 21453 6780 21465 6783
rect 21232 6752 21465 6780
rect 21232 6740 21238 6752
rect 21453 6749 21465 6752
rect 21499 6780 21511 6783
rect 21910 6780 21916 6792
rect 21499 6752 21916 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 20162 6644 20168 6656
rect 19904 6616 20168 6644
rect 20162 6604 20168 6616
rect 20220 6644 20226 6656
rect 20257 6647 20315 6653
rect 20257 6644 20269 6647
rect 20220 6616 20269 6644
rect 20220 6604 20226 6616
rect 20257 6613 20269 6616
rect 20303 6613 20315 6647
rect 21634 6644 21640 6656
rect 21595 6616 21640 6644
rect 20257 6607 20315 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 22060 6616 22293 6644
rect 22060 6604 22066 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 1104 6554 28336 6576
rect 1104 6502 1782 6554
rect 1834 6502 1846 6554
rect 1898 6502 1910 6554
rect 1962 6502 1974 6554
rect 2026 6502 4782 6554
rect 4834 6502 4846 6554
rect 4898 6502 4910 6554
rect 4962 6502 4974 6554
rect 5026 6502 7782 6554
rect 7834 6502 7846 6554
rect 7898 6502 7910 6554
rect 7962 6502 7974 6554
rect 8026 6502 10782 6554
rect 10834 6502 10846 6554
rect 10898 6502 10910 6554
rect 10962 6502 10974 6554
rect 11026 6502 13782 6554
rect 13834 6502 13846 6554
rect 13898 6502 13910 6554
rect 13962 6502 13974 6554
rect 14026 6502 16782 6554
rect 16834 6502 16846 6554
rect 16898 6502 16910 6554
rect 16962 6502 16974 6554
rect 17026 6502 19782 6554
rect 19834 6502 19846 6554
rect 19898 6502 19910 6554
rect 19962 6502 19974 6554
rect 20026 6502 22782 6554
rect 22834 6502 22846 6554
rect 22898 6502 22910 6554
rect 22962 6502 22974 6554
rect 23026 6502 25782 6554
rect 25834 6502 25846 6554
rect 25898 6502 25910 6554
rect 25962 6502 25974 6554
rect 26026 6502 28336 6554
rect 1104 6480 28336 6502
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 5368 6412 7205 6440
rect 5368 6384 5396 6412
rect 7193 6409 7205 6412
rect 7239 6440 7251 6443
rect 7466 6440 7472 6452
rect 7239 6412 7472 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 9582 6440 9588 6452
rect 9539 6412 9588 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 9582 6400 9588 6412
rect 9640 6440 9646 6452
rect 10042 6440 10048 6452
rect 9640 6412 10048 6440
rect 9640 6400 9646 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10652 6412 10701 6440
rect 10652 6400 10658 6412
rect 10689 6409 10701 6412
rect 10735 6440 10747 6443
rect 12158 6440 12164 6452
rect 10735 6412 12164 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 14093 6443 14151 6449
rect 14093 6440 14105 6443
rect 12768 6412 14105 6440
rect 12768 6400 12774 6412
rect 14093 6409 14105 6412
rect 14139 6440 14151 6443
rect 15838 6440 15844 6452
rect 14139 6412 15844 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 5350 6372 5356 6384
rect 5263 6344 5356 6372
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 5905 6375 5963 6381
rect 5905 6341 5917 6375
rect 5951 6372 5963 6375
rect 9769 6375 9827 6381
rect 5951 6344 8156 6372
rect 5951 6341 5963 6344
rect 5905 6335 5963 6341
rect 8128 6316 8156 6344
rect 9769 6341 9781 6375
rect 9815 6372 9827 6375
rect 9858 6372 9864 6384
rect 9815 6344 9864 6372
rect 9815 6341 9827 6344
rect 9769 6335 9827 6341
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 11057 6375 11115 6381
rect 11057 6341 11069 6375
rect 11103 6372 11115 6375
rect 11698 6372 11704 6384
rect 11103 6344 11704 6372
rect 11103 6341 11115 6344
rect 11057 6335 11115 6341
rect 11698 6332 11704 6344
rect 11756 6372 11762 6384
rect 12621 6375 12679 6381
rect 12621 6372 12633 6375
rect 11756 6344 12633 6372
rect 11756 6332 11762 6344
rect 12621 6341 12633 6344
rect 12667 6341 12679 6375
rect 12621 6335 12679 6341
rect 15289 6375 15347 6381
rect 15289 6341 15301 6375
rect 15335 6372 15347 6375
rect 15654 6372 15660 6384
rect 15335 6344 15660 6372
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 15654 6332 15660 6344
rect 15712 6332 15718 6384
rect 16117 6375 16175 6381
rect 16117 6341 16129 6375
rect 16163 6372 16175 6375
rect 18325 6375 18383 6381
rect 18325 6372 18337 6375
rect 16163 6344 18337 6372
rect 16163 6341 16175 6344
rect 16117 6335 16175 6341
rect 18325 6341 18337 6344
rect 18371 6372 18383 6375
rect 18874 6372 18880 6384
rect 18371 6344 18880 6372
rect 18371 6341 18383 6344
rect 18325 6335 18383 6341
rect 18874 6332 18880 6344
rect 18932 6372 18938 6384
rect 18932 6344 19380 6372
rect 18932 6332 18938 6344
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 6270 6304 6276 6316
rect 6231 6276 6276 6304
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 7650 6264 7656 6316
rect 7708 6304 7714 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7708 6276 7941 6304
rect 7708 6264 7714 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 8110 6304 8116 6316
rect 8023 6276 8116 6304
rect 7929 6267 7987 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 8294 6304 8300 6316
rect 8255 6276 8300 6304
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8754 6304 8760 6316
rect 8667 6276 8760 6304
rect 8754 6264 8760 6276
rect 8812 6304 8818 6316
rect 9950 6304 9956 6316
rect 8812 6276 8984 6304
rect 9911 6276 9956 6304
rect 8812 6264 8818 6276
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 7064 6208 7481 6236
rect 7064 6196 7070 6208
rect 7469 6205 7481 6208
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 8662 6196 8668 6248
rect 8720 6236 8726 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8720 6208 8861 6236
rect 8720 6196 8726 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8956 6236 8984 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 11330 6304 11336 6316
rect 11291 6276 11336 6304
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11790 6304 11796 6316
rect 11751 6276 11796 6304
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13446 6304 13452 6316
rect 13407 6276 13452 6304
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14366 6304 14372 6316
rect 14327 6276 14372 6304
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14461 6307 14519 6313
rect 14461 6273 14473 6307
rect 14507 6304 14519 6307
rect 14642 6304 14648 6316
rect 14507 6276 14648 6304
rect 14507 6273 14519 6276
rect 14461 6267 14519 6273
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 19352 6313 19380 6344
rect 21634 6332 21640 6384
rect 21692 6332 21698 6384
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 15988 6276 16957 6304
rect 15988 6264 15994 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 19518 6264 19524 6316
rect 19576 6304 19582 6316
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19576 6276 19717 6304
rect 19576 6264 19582 6276
rect 19705 6273 19717 6276
rect 19751 6304 19763 6307
rect 20622 6304 20628 6316
rect 19751 6276 20628 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 8956 6208 10241 6236
rect 8849 6199 8907 6205
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 13538 6236 13544 6248
rect 13499 6208 13544 6236
rect 10229 6199 10287 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16632 6208 16681 6236
rect 16632 6196 16638 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 17126 6236 17132 6248
rect 17087 6208 17132 6236
rect 16669 6199 16727 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6205 19487 6239
rect 19610 6236 19616 6248
rect 19523 6208 19616 6236
rect 19429 6199 19487 6205
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 8352 6140 11529 6168
rect 8352 6128 8358 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 11517 6131 11575 6137
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 19444 6168 19472 6199
rect 19610 6196 19616 6208
rect 19668 6236 19674 6248
rect 20165 6239 20223 6245
rect 20165 6236 20177 6239
rect 19668 6208 20177 6236
rect 19668 6196 19674 6208
rect 20165 6205 20177 6208
rect 20211 6205 20223 6239
rect 20714 6236 20720 6248
rect 20675 6208 20720 6236
rect 20165 6199 20223 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 20990 6236 20996 6248
rect 20951 6208 20996 6236
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22060 6208 22753 6236
rect 22060 6196 22066 6208
rect 22741 6205 22753 6208
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 20070 6168 20076 6180
rect 18840 6140 20076 6168
rect 18840 6128 18846 6140
rect 20070 6128 20076 6140
rect 20128 6128 20134 6180
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 14645 6103 14703 6109
rect 14645 6100 14657 6103
rect 14516 6072 14657 6100
rect 14516 6060 14522 6072
rect 14645 6069 14657 6072
rect 14691 6069 14703 6103
rect 14645 6063 14703 6069
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 16724 6072 17417 6100
rect 16724 6060 16730 6072
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 18966 6100 18972 6112
rect 18927 6072 18972 6100
rect 17405 6063 17463 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 1104 6010 28336 6032
rect 1104 5958 3282 6010
rect 3334 5958 3346 6010
rect 3398 5958 3410 6010
rect 3462 5958 3474 6010
rect 3526 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 6410 6010
rect 6462 5958 6474 6010
rect 6526 5958 9282 6010
rect 9334 5958 9346 6010
rect 9398 5958 9410 6010
rect 9462 5958 9474 6010
rect 9526 5958 12282 6010
rect 12334 5958 12346 6010
rect 12398 5958 12410 6010
rect 12462 5958 12474 6010
rect 12526 5958 15282 6010
rect 15334 5958 15346 6010
rect 15398 5958 15410 6010
rect 15462 5958 15474 6010
rect 15526 5958 18282 6010
rect 18334 5958 18346 6010
rect 18398 5958 18410 6010
rect 18462 5958 18474 6010
rect 18526 5958 21282 6010
rect 21334 5958 21346 6010
rect 21398 5958 21410 6010
rect 21462 5958 21474 6010
rect 21526 5958 24282 6010
rect 24334 5958 24346 6010
rect 24398 5958 24410 6010
rect 24462 5958 24474 6010
rect 24526 5958 27282 6010
rect 27334 5958 27346 6010
rect 27398 5958 27410 6010
rect 27462 5958 27474 6010
rect 27526 5958 28336 6010
rect 1104 5936 28336 5958
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5592 5868 5825 5896
rect 5592 5856 5598 5868
rect 5813 5865 5825 5868
rect 5859 5896 5871 5899
rect 6822 5896 6828 5908
rect 5859 5868 6828 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 7708 5868 9045 5896
rect 7708 5856 7714 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 10965 5899 11023 5905
rect 10965 5865 10977 5899
rect 11011 5896 11023 5899
rect 11330 5896 11336 5908
rect 11011 5868 11336 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 18509 5899 18567 5905
rect 14415 5868 18276 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 10597 5831 10655 5837
rect 10597 5797 10609 5831
rect 10643 5828 10655 5831
rect 12986 5828 12992 5840
rect 10643 5800 12992 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 17954 5828 17960 5840
rect 16684 5800 17960 5828
rect 6730 5760 6736 5772
rect 6691 5732 6736 5760
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7006 5760 7012 5772
rect 6967 5732 7012 5760
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5760 8815 5763
rect 9122 5760 9128 5772
rect 8803 5732 9128 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 11977 5763 12035 5769
rect 11977 5729 11989 5763
rect 12023 5760 12035 5763
rect 13078 5760 13084 5772
rect 12023 5732 13084 5760
rect 12023 5729 12035 5732
rect 11977 5723 12035 5729
rect 13078 5720 13084 5732
rect 13136 5760 13142 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13136 5732 13645 5760
rect 13136 5720 13142 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14458 5720 14464 5772
rect 14516 5760 14522 5772
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 14516 5732 16037 5760
rect 14516 5720 14522 5732
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16025 5723 16083 5729
rect 16206 5720 16212 5772
rect 16264 5760 16270 5772
rect 16577 5763 16635 5769
rect 16577 5760 16589 5763
rect 16264 5732 16589 5760
rect 16264 5720 16270 5732
rect 16577 5729 16589 5732
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 9950 5692 9956 5704
rect 9863 5664 9956 5692
rect 9950 5652 9956 5664
rect 10008 5692 10014 5704
rect 12802 5692 12808 5704
rect 10008 5664 11652 5692
rect 12763 5664 12808 5692
rect 10008 5652 10014 5664
rect 11624 5636 11652 5664
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 12986 5692 12992 5704
rect 12943 5664 12992 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 14185 5695 14243 5701
rect 14185 5661 14197 5695
rect 14231 5692 14243 5695
rect 14274 5692 14280 5704
rect 14231 5664 14280 5692
rect 14231 5661 14243 5664
rect 14185 5655 14243 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 15930 5652 15936 5704
rect 15988 5692 15994 5704
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15988 5664 16129 5692
rect 15988 5652 15994 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 16117 5655 16175 5661
rect 16482 5652 16488 5664
rect 16540 5692 16546 5704
rect 16684 5692 16712 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 18248 5828 18276 5868
rect 18509 5865 18521 5899
rect 18555 5896 18567 5899
rect 19518 5896 19524 5908
rect 18555 5868 19524 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20533 5899 20591 5905
rect 20533 5865 20545 5899
rect 20579 5896 20591 5899
rect 20714 5896 20720 5908
rect 20579 5868 20720 5896
rect 20579 5865 20591 5868
rect 20533 5859 20591 5865
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 21174 5828 21180 5840
rect 18248 5800 21180 5828
rect 21174 5788 21180 5800
rect 21232 5788 21238 5840
rect 18782 5760 18788 5772
rect 18743 5732 18788 5760
rect 18782 5720 18788 5732
rect 18840 5720 18846 5772
rect 20165 5763 20223 5769
rect 20165 5729 20177 5763
rect 20211 5760 20223 5763
rect 20990 5760 20996 5772
rect 20211 5732 20996 5760
rect 20211 5729 20223 5732
rect 20165 5723 20223 5729
rect 20990 5720 20996 5732
rect 21048 5760 21054 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 21048 5732 21097 5760
rect 21048 5720 21054 5732
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 21818 5760 21824 5772
rect 21779 5732 21824 5760
rect 21085 5723 21143 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 22002 5760 22008 5772
rect 21963 5732 22008 5760
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 16540 5664 16712 5692
rect 16540 5652 16546 5664
rect 17126 5652 17132 5704
rect 17184 5692 17190 5704
rect 17405 5695 17463 5701
rect 17405 5692 17417 5695
rect 17184 5664 17417 5692
rect 17184 5652 17190 5664
rect 17405 5661 17417 5664
rect 17451 5692 17463 5695
rect 17773 5695 17831 5701
rect 17773 5692 17785 5695
rect 17451 5664 17785 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 17773 5661 17785 5664
rect 17819 5692 17831 5695
rect 17954 5692 17960 5704
rect 17819 5664 17960 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 17954 5652 17960 5664
rect 18012 5692 18018 5704
rect 18598 5692 18604 5704
rect 18012 5664 18604 5692
rect 18012 5652 18018 5664
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 18932 5664 19625 5692
rect 18932 5652 18938 5664
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 21726 5692 21732 5704
rect 21687 5664 21732 5692
rect 19613 5655 19671 5661
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 22097 5695 22155 5701
rect 22097 5661 22109 5695
rect 22143 5661 22155 5695
rect 22097 5655 22155 5661
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 11238 5624 11244 5636
rect 6696 5596 7512 5624
rect 11199 5596 11244 5624
rect 6696 5584 6702 5596
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 11422 5624 11428 5636
rect 11383 5596 11428 5624
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 11606 5624 11612 5636
rect 11567 5596 11612 5624
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 13357 5627 13415 5633
rect 13357 5624 13369 5627
rect 11716 5596 13369 5624
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5556 6515 5559
rect 8662 5556 8668 5568
rect 6503 5528 8668 5556
rect 6503 5525 6515 5528
rect 6457 5519 6515 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 11716 5556 11744 5596
rect 13357 5593 13369 5596
rect 13403 5593 13415 5627
rect 13357 5587 13415 5593
rect 15473 5627 15531 5633
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 16022 5624 16028 5636
rect 15519 5596 16028 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 19337 5627 19395 5633
rect 19337 5593 19349 5627
rect 19383 5624 19395 5627
rect 21358 5624 21364 5636
rect 19383 5596 21364 5624
rect 19383 5593 19395 5596
rect 19337 5587 19395 5593
rect 21358 5584 21364 5596
rect 21416 5624 21422 5636
rect 22112 5624 22140 5655
rect 21416 5596 22140 5624
rect 21416 5584 21422 5596
rect 11572 5528 11744 5556
rect 12529 5559 12587 5565
rect 11572 5516 11578 5528
rect 12529 5525 12541 5559
rect 12575 5556 12587 5559
rect 13538 5556 13544 5568
rect 12575 5528 13544 5556
rect 12575 5525 12587 5528
rect 12529 5519 12587 5525
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 16632 5528 16957 5556
rect 16632 5516 16638 5528
rect 16945 5525 16957 5528
rect 16991 5525 17003 5559
rect 16945 5519 17003 5525
rect 1104 5466 28336 5488
rect 1104 5414 1782 5466
rect 1834 5414 1846 5466
rect 1898 5414 1910 5466
rect 1962 5414 1974 5466
rect 2026 5414 4782 5466
rect 4834 5414 4846 5466
rect 4898 5414 4910 5466
rect 4962 5414 4974 5466
rect 5026 5414 7782 5466
rect 7834 5414 7846 5466
rect 7898 5414 7910 5466
rect 7962 5414 7974 5466
rect 8026 5414 10782 5466
rect 10834 5414 10846 5466
rect 10898 5414 10910 5466
rect 10962 5414 10974 5466
rect 11026 5414 13782 5466
rect 13834 5414 13846 5466
rect 13898 5414 13910 5466
rect 13962 5414 13974 5466
rect 14026 5414 16782 5466
rect 16834 5414 16846 5466
rect 16898 5414 16910 5466
rect 16962 5414 16974 5466
rect 17026 5414 19782 5466
rect 19834 5414 19846 5466
rect 19898 5414 19910 5466
rect 19962 5414 19974 5466
rect 20026 5414 22782 5466
rect 22834 5414 22846 5466
rect 22898 5414 22910 5466
rect 22962 5414 22974 5466
rect 23026 5414 25782 5466
rect 25834 5414 25846 5466
rect 25898 5414 25910 5466
rect 25962 5414 25974 5466
rect 26026 5414 28336 5466
rect 1104 5392 28336 5414
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6638 5352 6644 5364
rect 6503 5324 6644 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7064 5324 7389 5352
rect 7064 5312 7070 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 8110 5352 8116 5364
rect 8071 5324 8116 5352
rect 7377 5315 7435 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 14277 5355 14335 5361
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 15930 5352 15936 5364
rect 14323 5324 15936 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 15930 5312 15936 5324
rect 15988 5352 15994 5364
rect 17313 5355 17371 5361
rect 17313 5352 17325 5355
rect 15988 5324 17325 5352
rect 15988 5312 15994 5324
rect 17313 5321 17325 5324
rect 17359 5321 17371 5355
rect 17313 5315 17371 5321
rect 18325 5355 18383 5361
rect 18325 5321 18337 5355
rect 18371 5352 18383 5355
rect 18598 5352 18604 5364
rect 18371 5324 18604 5352
rect 18371 5321 18383 5324
rect 18325 5315 18383 5321
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 21085 5355 21143 5361
rect 21085 5321 21097 5355
rect 21131 5352 21143 5355
rect 21634 5352 21640 5364
rect 21131 5324 21640 5352
rect 21131 5321 21143 5324
rect 21085 5315 21143 5321
rect 21634 5312 21640 5324
rect 21692 5312 21698 5364
rect 21818 5352 21824 5364
rect 21779 5324 21824 5352
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 7837 5287 7895 5293
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 8294 5284 8300 5296
rect 7883 5256 8300 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8662 5284 8668 5296
rect 8623 5256 8668 5284
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 11606 5284 11612 5296
rect 9180 5256 9720 5284
rect 11519 5256 11612 5284
rect 9180 5244 9186 5256
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7009 5219 7067 5225
rect 7009 5216 7021 5219
rect 6788 5188 7021 5216
rect 6788 5176 6794 5188
rect 7009 5185 7021 5188
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9582 5216 9588 5228
rect 9539 5188 9588 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 9692 5225 9720 5256
rect 11606 5244 11612 5256
rect 11664 5284 11670 5296
rect 14918 5284 14924 5296
rect 11664 5256 14924 5284
rect 11664 5244 11670 5256
rect 14918 5244 14924 5256
rect 14976 5244 14982 5296
rect 16666 5284 16672 5296
rect 16627 5256 16672 5284
rect 16666 5244 16672 5256
rect 16724 5244 16730 5296
rect 18966 5284 18972 5296
rect 18927 5256 18972 5284
rect 18966 5244 18972 5256
rect 19024 5244 19030 5296
rect 19702 5244 19708 5296
rect 19760 5244 19766 5296
rect 21358 5284 21364 5296
rect 21319 5256 21364 5284
rect 21358 5244 21364 5256
rect 21416 5244 21422 5296
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5185 9735 5219
rect 11146 5216 11152 5228
rect 11107 5188 11152 5216
rect 9677 5179 9735 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11422 5216 11428 5228
rect 11287 5188 11428 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11422 5176 11428 5188
rect 11480 5216 11486 5228
rect 11882 5216 11888 5228
rect 11480 5188 11888 5216
rect 11480 5176 11486 5188
rect 11882 5176 11888 5188
rect 11940 5216 11946 5228
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 11940 5188 12633 5216
rect 11940 5176 11946 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 12621 5179 12679 5185
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 14642 5216 14648 5228
rect 13403 5188 14648 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 15657 5219 15715 5225
rect 15657 5216 15669 5219
rect 15335 5188 15669 5216
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15657 5185 15669 5188
rect 15703 5216 15715 5219
rect 16206 5216 16212 5228
rect 16264 5225 16270 5228
rect 16264 5219 16287 5225
rect 15703 5188 16212 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 16206 5176 16212 5188
rect 16275 5216 16287 5219
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16275 5188 16957 5216
rect 16275 5185 16287 5188
rect 16264 5179 16287 5185
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 16264 5176 16270 5179
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 12710 5148 12716 5160
rect 12671 5120 12716 5148
rect 9217 5111 9275 5117
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 9232 5080 9260 5111
rect 12710 5108 12716 5120
rect 12768 5148 12774 5160
rect 12986 5148 12992 5160
rect 12768 5120 12992 5148
rect 12768 5108 12774 5120
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 16117 5151 16175 5157
rect 16117 5148 16129 5151
rect 14424 5120 16129 5148
rect 14424 5108 14430 5120
rect 16117 5117 16129 5120
rect 16163 5148 16175 5151
rect 17770 5148 17776 5160
rect 16163 5120 17776 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5148 18751 5151
rect 19058 5148 19064 5160
rect 18739 5120 19064 5148
rect 18739 5117 18751 5120
rect 18693 5111 18751 5117
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 20162 5108 20168 5160
rect 20220 5148 20226 5160
rect 20717 5151 20775 5157
rect 20717 5148 20729 5151
rect 20220 5120 20729 5148
rect 20220 5108 20226 5120
rect 20717 5117 20729 5120
rect 20763 5117 20775 5151
rect 20717 5111 20775 5117
rect 11238 5080 11244 5092
rect 9180 5052 11244 5080
rect 9180 5040 9186 5052
rect 11238 5040 11244 5052
rect 11296 5080 11302 5092
rect 11885 5083 11943 5089
rect 11885 5080 11897 5083
rect 11296 5052 11897 5080
rect 11296 5040 11302 5052
rect 11885 5049 11897 5052
rect 11931 5080 11943 5083
rect 18598 5080 18604 5092
rect 11931 5052 18604 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 10226 5012 10232 5024
rect 10187 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 14734 5012 14740 5024
rect 13955 4984 14740 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 14734 4972 14740 4984
rect 14792 5012 14798 5024
rect 16482 5012 16488 5024
rect 14792 4984 16488 5012
rect 14792 4972 14798 4984
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 1104 4922 28336 4944
rect 1104 4870 3282 4922
rect 3334 4870 3346 4922
rect 3398 4870 3410 4922
rect 3462 4870 3474 4922
rect 3526 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 6410 4922
rect 6462 4870 6474 4922
rect 6526 4870 9282 4922
rect 9334 4870 9346 4922
rect 9398 4870 9410 4922
rect 9462 4870 9474 4922
rect 9526 4870 12282 4922
rect 12334 4870 12346 4922
rect 12398 4870 12410 4922
rect 12462 4870 12474 4922
rect 12526 4870 15282 4922
rect 15334 4870 15346 4922
rect 15398 4870 15410 4922
rect 15462 4870 15474 4922
rect 15526 4870 18282 4922
rect 18334 4870 18346 4922
rect 18398 4870 18410 4922
rect 18462 4870 18474 4922
rect 18526 4870 21282 4922
rect 21334 4870 21346 4922
rect 21398 4870 21410 4922
rect 21462 4870 21474 4922
rect 21526 4870 24282 4922
rect 24334 4870 24346 4922
rect 24398 4870 24410 4922
rect 24462 4870 24474 4922
rect 24526 4870 27282 4922
rect 27334 4870 27346 4922
rect 27398 4870 27410 4922
rect 27462 4870 27474 4922
rect 27526 4870 28336 4922
rect 1104 4848 28336 4870
rect 6822 4808 6828 4820
rect 6783 4780 6828 4808
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 8754 4808 8760 4820
rect 7607 4780 8760 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9122 4808 9128 4820
rect 9083 4780 9128 4808
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 11882 4808 11888 4820
rect 11843 4780 11888 4808
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 13909 4811 13967 4817
rect 13909 4777 13921 4811
rect 13955 4808 13967 4811
rect 14458 4808 14464 4820
rect 13955 4780 14464 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 18325 4811 18383 4817
rect 18325 4777 18337 4811
rect 18371 4808 18383 4811
rect 18966 4808 18972 4820
rect 18371 4780 18972 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19702 4768 19708 4820
rect 19760 4808 19766 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19760 4780 19809 4808
rect 19760 4768 19766 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 20162 4808 20168 4820
rect 20123 4780 20168 4808
rect 19797 4771 19855 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 21545 4811 21603 4817
rect 21545 4777 21557 4811
rect 21591 4808 21603 4811
rect 22002 4808 22008 4820
rect 21591 4780 22008 4808
rect 21591 4777 21603 4780
rect 21545 4771 21603 4777
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 18598 4700 18604 4752
rect 18656 4740 18662 4752
rect 18785 4743 18843 4749
rect 18785 4740 18797 4743
rect 18656 4712 18797 4740
rect 18656 4700 18662 4712
rect 18785 4709 18797 4712
rect 18831 4709 18843 4743
rect 18785 4703 18843 4709
rect 19058 4700 19064 4752
rect 19116 4740 19122 4752
rect 19153 4743 19211 4749
rect 19153 4740 19165 4743
rect 19116 4712 19165 4740
rect 19116 4700 19122 4712
rect 19153 4709 19165 4712
rect 19199 4740 19211 4743
rect 20714 4740 20720 4752
rect 19199 4712 20720 4740
rect 19199 4709 19211 4712
rect 19153 4703 19211 4709
rect 20714 4700 20720 4712
rect 20772 4700 20778 4752
rect 21177 4743 21235 4749
rect 21177 4709 21189 4743
rect 21223 4740 21235 4743
rect 21726 4740 21732 4752
rect 21223 4712 21732 4740
rect 21223 4709 21235 4712
rect 21177 4703 21235 4709
rect 21726 4700 21732 4712
rect 21784 4700 21790 4752
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 10042 4672 10048 4684
rect 7975 4644 9628 4672
rect 9955 4644 10048 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 9600 4616 9628 4644
rect 10042 4632 10048 4644
rect 10100 4672 10106 4684
rect 14001 4675 14059 4681
rect 10100 4644 11376 4672
rect 10100 4632 10106 4644
rect 8294 4604 8300 4616
rect 7116 4576 8300 4604
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 7116 4477 7144 4576
rect 8294 4564 8300 4576
rect 8352 4613 8358 4616
rect 8352 4607 8407 4613
rect 8352 4573 8361 4607
rect 8395 4573 8407 4607
rect 8352 4567 8407 4573
rect 8352 4564 8358 4567
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 9640 4576 10333 4604
rect 9640 4564 9646 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10321 4567 10379 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11146 4604 11152 4616
rect 11011 4576 11152 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 8205 4539 8263 4545
rect 8205 4536 8217 4539
rect 8168 4508 8217 4536
rect 8168 4496 8174 4508
rect 8205 4505 8217 4508
rect 8251 4505 8263 4539
rect 8205 4499 8263 4505
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10796 4536 10824 4567
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11348 4613 11376 4644
rect 14001 4641 14013 4675
rect 14047 4672 14059 4675
rect 14274 4672 14280 4684
rect 14047 4644 14280 4672
rect 14047 4641 14059 4644
rect 14001 4635 14059 4641
rect 14274 4632 14280 4644
rect 14332 4672 14338 4684
rect 15010 4672 15016 4684
rect 14332 4644 15016 4672
rect 14332 4632 14338 4644
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 16022 4672 16028 4684
rect 15983 4644 16028 4672
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 17770 4672 17776 4684
rect 17731 4644 17776 4672
rect 17770 4632 17776 4644
rect 17828 4632 17834 4684
rect 18138 4632 18144 4684
rect 18196 4672 18202 4684
rect 18874 4672 18880 4684
rect 18196 4644 18880 4672
rect 18196 4632 18202 4644
rect 18874 4632 18880 4644
rect 18932 4672 18938 4684
rect 18932 4644 19656 4672
rect 18932 4632 18938 4644
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 11422 4604 11428 4616
rect 11379 4576 11428 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 11882 4604 11888 4616
rect 11563 4576 11888 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 12066 4604 12072 4616
rect 11979 4576 12072 4604
rect 11992 4536 12020 4576
rect 12066 4564 12072 4576
rect 12124 4604 12130 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 12124 4576 13001 4604
rect 12124 4564 12130 4576
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 13170 4604 13176 4616
rect 13035 4576 13176 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 14194 4607 14252 4613
rect 14194 4573 14206 4607
rect 14240 4604 14252 4607
rect 14366 4604 14372 4616
rect 14240 4576 14372 4604
rect 14240 4573 14252 4576
rect 14194 4567 14252 4573
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 9548 4508 10456 4536
rect 10796 4508 12020 4536
rect 9548 4496 9554 4508
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 6696 4440 7113 4468
rect 6696 4428 6702 4440
rect 7101 4437 7113 4440
rect 7147 4437 7159 4471
rect 8478 4468 8484 4480
rect 8439 4440 8484 4468
rect 7101 4431 7159 4437
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 10428 4468 10456 4508
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 13081 4539 13139 4545
rect 13081 4536 13093 4539
rect 12768 4508 13093 4536
rect 12768 4496 12774 4508
rect 13081 4505 13093 4508
rect 13127 4536 13139 4539
rect 13354 4536 13360 4548
rect 13127 4508 13360 4536
rect 13127 4505 13139 4508
rect 13081 4499 13139 4505
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 13541 4539 13599 4545
rect 13541 4505 13553 4539
rect 13587 4536 13599 4539
rect 14001 4539 14059 4545
rect 14001 4536 14013 4539
rect 13587 4508 14013 4536
rect 13587 4505 13599 4508
rect 13541 4499 13599 4505
rect 14001 4505 14013 4508
rect 14047 4505 14059 4539
rect 14001 4499 14059 4505
rect 15764 4480 15792 4567
rect 17126 4564 17132 4616
rect 17184 4564 17190 4616
rect 18598 4604 18604 4616
rect 18559 4576 18604 4604
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 19628 4613 19656 4644
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 11146 4468 11152 4480
rect 10428 4440 11152 4468
rect 11146 4428 11152 4440
rect 11204 4468 11210 4480
rect 12986 4468 12992 4480
rect 11204 4440 12992 4468
rect 11204 4428 11210 4440
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 14369 4471 14427 4477
rect 14369 4468 14381 4471
rect 13688 4440 14381 4468
rect 13688 4428 13694 4440
rect 14369 4437 14381 4440
rect 14415 4437 14427 4471
rect 15746 4468 15752 4480
rect 15659 4440 15752 4468
rect 14369 4431 14427 4437
rect 15746 4428 15752 4440
rect 15804 4468 15810 4480
rect 19058 4468 19064 4480
rect 15804 4440 19064 4468
rect 15804 4428 15810 4440
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 20162 4428 20168 4480
rect 20220 4468 20226 4480
rect 20441 4471 20499 4477
rect 20441 4468 20453 4471
rect 20220 4440 20453 4468
rect 20220 4428 20226 4440
rect 20441 4437 20453 4440
rect 20487 4437 20499 4471
rect 20441 4431 20499 4437
rect 1104 4378 28336 4400
rect 1104 4326 1782 4378
rect 1834 4326 1846 4378
rect 1898 4326 1910 4378
rect 1962 4326 1974 4378
rect 2026 4326 4782 4378
rect 4834 4326 4846 4378
rect 4898 4326 4910 4378
rect 4962 4326 4974 4378
rect 5026 4326 7782 4378
rect 7834 4326 7846 4378
rect 7898 4326 7910 4378
rect 7962 4326 7974 4378
rect 8026 4326 10782 4378
rect 10834 4326 10846 4378
rect 10898 4326 10910 4378
rect 10962 4326 10974 4378
rect 11026 4326 13782 4378
rect 13834 4326 13846 4378
rect 13898 4326 13910 4378
rect 13962 4326 13974 4378
rect 14026 4326 16782 4378
rect 16834 4326 16846 4378
rect 16898 4326 16910 4378
rect 16962 4326 16974 4378
rect 17026 4326 19782 4378
rect 19834 4326 19846 4378
rect 19898 4326 19910 4378
rect 19962 4326 19974 4378
rect 20026 4326 22782 4378
rect 22834 4326 22846 4378
rect 22898 4326 22910 4378
rect 22962 4326 22974 4378
rect 23026 4326 25782 4378
rect 25834 4326 25846 4378
rect 25898 4326 25910 4378
rect 25962 4326 25974 4378
rect 26026 4326 28336 4378
rect 1104 4304 28336 4326
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11882 4264 11888 4276
rect 10735 4236 11888 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 11882 4224 11888 4236
rect 11940 4264 11946 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11940 4236 11989 4264
rect 11940 4224 11946 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 11977 4227 12035 4233
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 14921 4267 14979 4273
rect 14921 4264 14933 4267
rect 13596 4236 14933 4264
rect 13596 4224 13602 4236
rect 14921 4233 14933 4236
rect 14967 4233 14979 4267
rect 14921 4227 14979 4233
rect 15473 4267 15531 4273
rect 15473 4233 15485 4267
rect 15519 4264 15531 4267
rect 16022 4264 16028 4276
rect 15519 4236 16028 4264
rect 15519 4233 15531 4236
rect 15473 4227 15531 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 16298 4224 16304 4276
rect 16356 4264 16362 4276
rect 18693 4267 18751 4273
rect 18693 4264 18705 4267
rect 16356 4236 18705 4264
rect 16356 4224 16362 4236
rect 18693 4233 18705 4236
rect 18739 4233 18751 4267
rect 18693 4227 18751 4233
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19610 4264 19616 4276
rect 19383 4236 19616 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 8846 4196 8852 4208
rect 6788 4168 8852 4196
rect 6788 4156 6794 4168
rect 7650 4128 7656 4140
rect 7611 4100 7656 4128
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8312 4137 8340 4168
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 9030 4156 9036 4208
rect 9088 4156 9094 4208
rect 10226 4156 10232 4208
rect 10284 4196 10290 4208
rect 11609 4199 11667 4205
rect 11609 4196 11621 4199
rect 10284 4168 11621 4196
rect 10284 4156 10290 4168
rect 11609 4165 11621 4168
rect 11655 4196 11667 4199
rect 11790 4196 11796 4208
rect 11655 4168 11796 4196
rect 11655 4165 11667 4168
rect 11609 4159 11667 4165
rect 11790 4156 11796 4168
rect 11848 4196 11854 4208
rect 12713 4199 12771 4205
rect 12713 4196 12725 4199
rect 11848 4168 12725 4196
rect 11848 4156 11854 4168
rect 12713 4165 12725 4168
rect 12759 4196 12771 4199
rect 12894 4196 12900 4208
rect 12759 4168 12900 4196
rect 12759 4165 12771 4168
rect 12713 4159 12771 4165
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 12986 4156 12992 4208
rect 13044 4196 13050 4208
rect 14277 4199 14335 4205
rect 14277 4196 14289 4199
rect 13044 4168 14289 4196
rect 13044 4156 13050 4168
rect 14277 4165 14289 4168
rect 14323 4196 14335 4199
rect 16850 4196 16856 4208
rect 14323 4168 16856 4196
rect 14323 4165 14335 4168
rect 14277 4159 14335 4165
rect 16850 4156 16856 4168
rect 16908 4156 16914 4208
rect 18598 4196 18604 4208
rect 17512 4168 18604 4196
rect 17512 4140 17540 4168
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8275 4100 8309 4128
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 12805 4131 12863 4137
rect 12805 4128 12817 4131
rect 11204 4100 12817 4128
rect 11204 4088 11210 4100
rect 12805 4097 12817 4100
rect 12851 4128 12863 4131
rect 14001 4131 14059 4137
rect 12851 4100 13492 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 8570 4060 8576 4072
rect 8531 4032 8576 4060
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4029 10379 4063
rect 10321 4023 10379 4029
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 12710 4060 12716 4072
rect 11379 4032 12716 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6638 3924 6644 3936
rect 6503 3896 6644 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 8018 3924 8024 3936
rect 7979 3896 8024 3924
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9582 3924 9588 3936
rect 8352 3896 9588 3924
rect 8352 3884 8358 3896
rect 9582 3884 9588 3896
rect 9640 3924 9646 3936
rect 10336 3924 10364 4023
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 13464 4060 13492 4100
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14366 4128 14372 4140
rect 14047 4100 14372 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 16761 4131 16819 4137
rect 16761 4097 16773 4131
rect 16807 4128 16819 4131
rect 17494 4128 17500 4140
rect 16807 4100 17500 4128
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17954 4088 17960 4140
rect 18012 4128 18018 4140
rect 18524 4137 18552 4168
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 18233 4131 18291 4137
rect 18233 4128 18245 4131
rect 18012 4100 18245 4128
rect 18012 4088 18018 4100
rect 18233 4097 18245 4100
rect 18279 4097 18291 4131
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 18487 4100 18521 4128
rect 18233 4091 18291 4097
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 19610 4128 19616 4140
rect 18932 4100 19616 4128
rect 18932 4088 18938 4100
rect 19610 4088 19616 4100
rect 19668 4128 19674 4140
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19668 4100 20085 4128
rect 19668 4088 19674 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 13464 4032 14657 4060
rect 14645 4029 14657 4032
rect 14691 4060 14703 4063
rect 14918 4060 14924 4072
rect 14691 4032 14924 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 14918 4020 14924 4032
rect 14976 4060 14982 4072
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 14976 4032 17601 4060
rect 14976 4020 14982 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 17828 4032 18368 4060
rect 17828 4020 17834 4032
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 14458 4001 14464 4004
rect 14442 3995 14464 4001
rect 14442 3992 14454 3995
rect 13228 3964 14044 3992
rect 14371 3964 14454 3992
rect 13228 3952 13234 3964
rect 9640 3896 10364 3924
rect 14016 3924 14044 3964
rect 14442 3961 14454 3964
rect 14516 3992 14522 4004
rect 16574 3992 16580 4004
rect 14516 3964 16580 3992
rect 14442 3955 14464 3961
rect 14458 3952 14464 3955
rect 14516 3952 14522 3964
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 18340 4001 18368 4032
rect 17221 3995 17279 4001
rect 17221 3992 17233 3995
rect 17184 3964 17233 3992
rect 17184 3952 17190 3964
rect 17221 3961 17233 3964
rect 17267 3992 17279 3995
rect 18325 3995 18383 4001
rect 17267 3964 18276 3992
rect 17267 3961 17279 3964
rect 17221 3955 17279 3961
rect 14550 3924 14556 3936
rect 14016 3896 14556 3924
rect 9640 3884 9646 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 15746 3924 15752 3936
rect 15707 3896 15752 3924
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 18248 3924 18276 3964
rect 18325 3961 18337 3995
rect 18371 3992 18383 3995
rect 19334 3992 19340 4004
rect 18371 3964 19340 3992
rect 18371 3961 18383 3964
rect 18325 3955 18383 3961
rect 19334 3952 19340 3964
rect 19392 3952 19398 4004
rect 19797 3927 19855 3933
rect 19797 3924 19809 3927
rect 18248 3896 19809 3924
rect 19797 3893 19809 3896
rect 19843 3893 19855 3927
rect 20438 3924 20444 3936
rect 20399 3896 20444 3924
rect 19797 3887 19855 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 1104 3834 28336 3856
rect 1104 3782 3282 3834
rect 3334 3782 3346 3834
rect 3398 3782 3410 3834
rect 3462 3782 3474 3834
rect 3526 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 6410 3834
rect 6462 3782 6474 3834
rect 6526 3782 9282 3834
rect 9334 3782 9346 3834
rect 9398 3782 9410 3834
rect 9462 3782 9474 3834
rect 9526 3782 12282 3834
rect 12334 3782 12346 3834
rect 12398 3782 12410 3834
rect 12462 3782 12474 3834
rect 12526 3782 15282 3834
rect 15334 3782 15346 3834
rect 15398 3782 15410 3834
rect 15462 3782 15474 3834
rect 15526 3782 18282 3834
rect 18334 3782 18346 3834
rect 18398 3782 18410 3834
rect 18462 3782 18474 3834
rect 18526 3782 21282 3834
rect 21334 3782 21346 3834
rect 21398 3782 21410 3834
rect 21462 3782 21474 3834
rect 21526 3782 24282 3834
rect 24334 3782 24346 3834
rect 24398 3782 24410 3834
rect 24462 3782 24474 3834
rect 24526 3782 27282 3834
rect 27334 3782 27346 3834
rect 27398 3782 27410 3834
rect 27462 3782 27474 3834
rect 27526 3782 28336 3834
rect 1104 3760 28336 3782
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 7190 3720 7196 3732
rect 7055 3692 7196 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 7190 3680 7196 3692
rect 7248 3720 7254 3732
rect 11422 3720 11428 3732
rect 7248 3692 11428 3720
rect 7248 3680 7254 3692
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11790 3720 11796 3732
rect 11751 3692 11796 3720
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 14090 3720 14096 3732
rect 12952 3692 14096 3720
rect 12952 3680 12958 3692
rect 14090 3680 14096 3692
rect 14148 3720 14154 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14148 3692 14657 3720
rect 14148 3680 14154 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18012 3692 18153 3720
rect 18012 3680 18018 3692
rect 18141 3689 18153 3692
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 20073 3723 20131 3729
rect 20073 3720 20085 3723
rect 19392 3692 20085 3720
rect 19392 3680 19398 3692
rect 20073 3689 20085 3692
rect 20119 3720 20131 3723
rect 20162 3720 20168 3732
rect 20119 3692 20168 3720
rect 20119 3689 20131 3692
rect 20073 3683 20131 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 8076 3624 8708 3652
rect 8076 3612 8082 3624
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 7708 3556 7757 3584
rect 7708 3544 7714 3556
rect 7745 3553 7757 3556
rect 7791 3584 7803 3587
rect 8478 3584 8484 3596
rect 7791 3556 8484 3584
rect 7791 3553 7803 3556
rect 7745 3547 7803 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 8680 3593 8708 3624
rect 11330 3612 11336 3664
rect 11388 3652 11394 3664
rect 14369 3655 14427 3661
rect 14369 3652 14381 3655
rect 11388 3624 14381 3652
rect 11388 3612 11394 3624
rect 14369 3621 14381 3624
rect 14415 3652 14427 3655
rect 14458 3652 14464 3664
rect 14415 3624 14464 3652
rect 14415 3621 14427 3624
rect 14369 3615 14427 3621
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 16850 3612 16856 3664
rect 16908 3652 16914 3664
rect 19153 3655 19211 3661
rect 19153 3652 19165 3655
rect 16908 3624 19165 3652
rect 16908 3612 16914 3624
rect 19153 3621 19165 3624
rect 19199 3621 19211 3655
rect 19153 3615 19211 3621
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 8711 3556 10149 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 10137 3553 10149 3556
rect 10183 3584 10195 3587
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10183 3556 10977 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10965 3553 10977 3556
rect 11011 3584 11023 3587
rect 11011 3556 11376 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8352 3488 8585 3516
rect 8352 3476 8358 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 11238 3516 11244 3528
rect 11199 3488 11244 3516
rect 8573 3479 8631 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11348 3516 11376 3556
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 14274 3584 14280 3596
rect 11480 3556 11525 3584
rect 12084 3556 14280 3584
rect 11480 3544 11486 3556
rect 12084 3516 12112 3556
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 17494 3584 17500 3596
rect 17455 3556 17500 3584
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 11348 3488 12112 3516
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 7837 3451 7895 3457
rect 7837 3417 7849 3451
rect 7883 3448 7895 3451
rect 8478 3448 8484 3460
rect 7883 3420 8484 3448
rect 7883 3417 7895 3420
rect 7837 3411 7895 3417
rect 8478 3408 8484 3420
rect 8536 3408 8542 3460
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 9824 3420 10425 3448
rect 9824 3408 9830 3420
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 11256 3448 11284 3476
rect 12161 3451 12219 3457
rect 12161 3448 12173 3451
rect 11256 3420 12173 3448
rect 10413 3411 10471 3417
rect 12161 3417 12173 3420
rect 12207 3448 12219 3451
rect 12544 3448 12572 3479
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12952 3488 13093 3516
rect 12952 3476 12958 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 15746 3516 15752 3528
rect 13587 3488 13814 3516
rect 15707 3488 15752 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 12207 3420 12572 3448
rect 12207 3417 12219 3420
rect 12161 3411 12219 3417
rect 7374 3380 7380 3392
rect 7335 3352 7380 3380
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 8904 3352 9137 3380
rect 8904 3340 8910 3352
rect 9125 3349 9137 3352
rect 9171 3380 9183 3383
rect 9490 3380 9496 3392
rect 9171 3352 9496 3380
rect 9171 3349 9183 3352
rect 9125 3343 9183 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 13786 3380 13814 3488
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 16114 3516 16120 3528
rect 16075 3488 16120 3516
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 18690 3516 18696 3528
rect 18651 3488 18696 3516
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 17126 3408 17132 3460
rect 17184 3408 17190 3460
rect 14001 3383 14059 3389
rect 14001 3380 14013 3383
rect 13786 3352 14013 3380
rect 14001 3349 14013 3352
rect 14047 3380 14059 3383
rect 14182 3380 14188 3392
rect 14047 3352 14188 3380
rect 14047 3349 14059 3352
rect 14001 3343 14059 3349
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 18877 3383 18935 3389
rect 18877 3380 18889 3383
rect 18012 3352 18889 3380
rect 18012 3340 18018 3352
rect 18877 3349 18889 3352
rect 18923 3380 18935 3383
rect 19610 3380 19616 3392
rect 18923 3352 19616 3380
rect 18923 3349 18935 3352
rect 18877 3343 18935 3349
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 1104 3290 28336 3312
rect 1104 3238 1782 3290
rect 1834 3238 1846 3290
rect 1898 3238 1910 3290
rect 1962 3238 1974 3290
rect 2026 3238 4782 3290
rect 4834 3238 4846 3290
rect 4898 3238 4910 3290
rect 4962 3238 4974 3290
rect 5026 3238 7782 3290
rect 7834 3238 7846 3290
rect 7898 3238 7910 3290
rect 7962 3238 7974 3290
rect 8026 3238 10782 3290
rect 10834 3238 10846 3290
rect 10898 3238 10910 3290
rect 10962 3238 10974 3290
rect 11026 3238 13782 3290
rect 13834 3238 13846 3290
rect 13898 3238 13910 3290
rect 13962 3238 13974 3290
rect 14026 3238 16782 3290
rect 16834 3238 16846 3290
rect 16898 3238 16910 3290
rect 16962 3238 16974 3290
rect 17026 3238 19782 3290
rect 19834 3238 19846 3290
rect 19898 3238 19910 3290
rect 19962 3238 19974 3290
rect 20026 3238 22782 3290
rect 22834 3238 22846 3290
rect 22898 3238 22910 3290
rect 22962 3238 22974 3290
rect 23026 3238 25782 3290
rect 25834 3238 25846 3290
rect 25898 3238 25910 3290
rect 25962 3238 25974 3290
rect 26026 3238 28336 3290
rect 1104 3216 28336 3238
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3176 6515 3179
rect 6638 3176 6644 3188
rect 6503 3148 6644 3176
rect 6503 3145 6515 3148
rect 6457 3139 6515 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7469 3179 7527 3185
rect 7469 3145 7481 3179
rect 7515 3145 7527 3179
rect 7469 3139 7527 3145
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8110 3176 8116 3188
rect 7883 3148 8116 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 7484 3108 7512 3139
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 8570 3176 8576 3188
rect 8435 3148 8576 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9030 3176 9036 3188
rect 8803 3148 9036 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8772 3108 8800 3139
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 11422 3136 11428 3188
rect 11480 3176 11486 3188
rect 13078 3176 13084 3188
rect 11480 3148 13084 3176
rect 11480 3136 11486 3148
rect 9766 3108 9772 3120
rect 7484 3080 8800 3108
rect 9727 3080 9772 3108
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 10226 3068 10232 3120
rect 10284 3068 10290 3120
rect 11532 3117 11560 3148
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 16114 3176 16120 3188
rect 15519 3148 16120 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 19153 3179 19211 3185
rect 19153 3176 19165 3179
rect 18656 3148 19165 3176
rect 18656 3136 18662 3148
rect 19153 3145 19165 3148
rect 19199 3176 19211 3179
rect 19521 3179 19579 3185
rect 19521 3176 19533 3179
rect 19199 3148 19533 3176
rect 19199 3145 19211 3148
rect 19153 3139 19211 3145
rect 19521 3145 19533 3148
rect 19567 3176 19579 3179
rect 20438 3176 20444 3188
rect 19567 3148 20444 3176
rect 19567 3145 19579 3148
rect 19521 3139 19579 3145
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 11517 3111 11575 3117
rect 11517 3077 11529 3111
rect 11563 3077 11575 3111
rect 11517 3071 11575 3077
rect 12618 3068 12624 3120
rect 12676 3108 12682 3120
rect 13173 3111 13231 3117
rect 13173 3108 13185 3111
rect 12676 3080 13185 3108
rect 12676 3068 12682 3080
rect 13173 3077 13185 3080
rect 13219 3108 13231 3111
rect 13262 3108 13268 3120
rect 13219 3080 13268 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 13630 3068 13636 3120
rect 13688 3068 13694 3120
rect 14918 3108 14924 3120
rect 14879 3080 14924 3108
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 15010 3068 15016 3120
rect 15068 3108 15074 3120
rect 16393 3111 16451 3117
rect 16393 3108 16405 3111
rect 15068 3080 16405 3108
rect 15068 3068 15074 3080
rect 16393 3077 16405 3080
rect 16439 3108 16451 3111
rect 18690 3108 18696 3120
rect 16439 3080 18696 3108
rect 16439 3077 16451 3080
rect 16393 3071 16451 3077
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7374 3000 7380 3052
rect 7432 3040 7438 3052
rect 9122 3040 9128 3052
rect 7432 3012 9128 3040
rect 7432 3000 7438 3012
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 16942 3040 16948 3052
rect 16903 3012 16948 3040
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18012 3012 18245 3040
rect 18012 3000 18018 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 9490 2972 9496 2984
rect 9451 2944 9496 2972
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 12894 2972 12900 2984
rect 12807 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2972 12958 2984
rect 15746 2972 15752 2984
rect 12952 2944 15752 2972
rect 12952 2932 12958 2944
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 14424 2876 18429 2904
rect 14424 2864 14430 2876
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 18417 2867 18475 2873
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 13814 2836 13820 2848
rect 12115 2808 13820 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 13814 2796 13820 2808
rect 13872 2836 13878 2848
rect 14182 2836 14188 2848
rect 13872 2808 14188 2836
rect 13872 2796 13878 2808
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 17126 2796 17132 2848
rect 17184 2836 17190 2848
rect 17494 2836 17500 2848
rect 17184 2808 17500 2836
rect 17184 2796 17190 2808
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 1104 2746 28336 2768
rect 1104 2694 3282 2746
rect 3334 2694 3346 2746
rect 3398 2694 3410 2746
rect 3462 2694 3474 2746
rect 3526 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 6410 2746
rect 6462 2694 6474 2746
rect 6526 2694 9282 2746
rect 9334 2694 9346 2746
rect 9398 2694 9410 2746
rect 9462 2694 9474 2746
rect 9526 2694 12282 2746
rect 12334 2694 12346 2746
rect 12398 2694 12410 2746
rect 12462 2694 12474 2746
rect 12526 2694 15282 2746
rect 15334 2694 15346 2746
rect 15398 2694 15410 2746
rect 15462 2694 15474 2746
rect 15526 2694 18282 2746
rect 18334 2694 18346 2746
rect 18398 2694 18410 2746
rect 18462 2694 18474 2746
rect 18526 2694 21282 2746
rect 21334 2694 21346 2746
rect 21398 2694 21410 2746
rect 21462 2694 21474 2746
rect 21526 2694 24282 2746
rect 24334 2694 24346 2746
rect 24398 2694 24410 2746
rect 24462 2694 24474 2746
rect 24526 2694 27282 2746
rect 27334 2694 27346 2746
rect 27398 2694 27410 2746
rect 27462 2694 27474 2746
rect 27526 2694 28336 2746
rect 1104 2672 28336 2694
rect 7650 2632 7656 2644
rect 7611 2604 7656 2632
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9766 2632 9772 2644
rect 9079 2604 9772 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10226 2632 10232 2644
rect 10183 2604 10232 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 8665 2567 8723 2573
rect 8665 2533 8677 2567
rect 8711 2564 8723 2567
rect 10152 2564 10180 2595
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 11238 2632 11244 2644
rect 10551 2604 11244 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 11238 2592 11244 2604
rect 11296 2632 11302 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11296 2604 11437 2632
rect 11296 2592 11302 2604
rect 11425 2601 11437 2604
rect 11471 2601 11483 2635
rect 12894 2632 12900 2644
rect 12855 2604 12900 2632
rect 11425 2595 11483 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13262 2632 13268 2644
rect 13223 2604 13268 2632
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 17037 2635 17095 2641
rect 17037 2632 17049 2635
rect 13412 2604 17049 2632
rect 13412 2592 13418 2604
rect 8711 2536 10180 2564
rect 12253 2567 12311 2573
rect 8711 2533 8723 2536
rect 8665 2527 8723 2533
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 13630 2564 13636 2576
rect 12299 2536 13636 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 13924 2573 13952 2604
rect 17037 2601 17049 2604
rect 17083 2601 17095 2635
rect 17037 2595 17095 2601
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 18877 2635 18935 2641
rect 18877 2632 18889 2635
rect 17552 2604 18889 2632
rect 17552 2592 17558 2604
rect 18877 2601 18889 2604
rect 18923 2601 18935 2635
rect 18877 2595 18935 2601
rect 13909 2567 13967 2573
rect 13909 2533 13921 2567
rect 13955 2533 13967 2567
rect 13909 2527 13967 2533
rect 14550 2524 14556 2576
rect 14608 2564 14614 2576
rect 17405 2567 17463 2573
rect 17405 2564 17417 2567
rect 14608 2536 17417 2564
rect 14608 2524 14614 2536
rect 17405 2533 17417 2536
rect 17451 2533 17463 2567
rect 17954 2564 17960 2576
rect 17915 2536 17960 2564
rect 17405 2527 17463 2533
rect 17954 2524 17960 2536
rect 18012 2524 18018 2576
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2496 10931 2499
rect 10919 2468 15148 2496
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7340 2400 7389 2428
rect 7340 2388 7346 2400
rect 7377 2397 7389 2400
rect 7423 2428 7435 2431
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 7423 2400 8309 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 8297 2397 8309 2400
rect 8343 2428 8355 2431
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 8343 2400 9965 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 9953 2397 9965 2400
rect 9999 2428 10011 2431
rect 10042 2428 10048 2440
rect 9999 2400 10048 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 11146 2428 11152 2440
rect 11059 2400 11152 2428
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 11256 2437 11284 2468
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14090 2428 14096 2440
rect 13872 2400 13965 2428
rect 14051 2400 14096 2428
rect 13872 2388 13878 2400
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 15120 2437 15148 2468
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 16298 2428 16304 2440
rect 15151 2400 16304 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 17972 2428 18000 2524
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 17972 2400 18705 2428
rect 18693 2397 18705 2400
rect 18739 2428 18751 2431
rect 19153 2431 19211 2437
rect 19153 2428 19165 2431
rect 18739 2400 19165 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 19153 2397 19165 2400
rect 19199 2397 19211 2431
rect 19153 2391 19211 2397
rect 9122 2320 9128 2372
rect 9180 2360 9186 2372
rect 11164 2360 11192 2388
rect 9180 2332 11192 2360
rect 13832 2360 13860 2388
rect 15657 2363 15715 2369
rect 15657 2360 15669 2363
rect 13832 2332 15669 2360
rect 9180 2320 9186 2332
rect 15657 2329 15669 2332
rect 15703 2329 15715 2363
rect 15657 2323 15715 2329
rect 16761 2363 16819 2369
rect 16761 2329 16773 2363
rect 16807 2360 16819 2363
rect 16942 2360 16948 2372
rect 16807 2332 16948 2360
rect 16807 2329 16819 2332
rect 16761 2323 16819 2329
rect 16942 2320 16948 2332
rect 17000 2360 17006 2372
rect 18230 2360 18236 2372
rect 17000 2332 18236 2360
rect 17000 2320 17006 2332
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2292 9370 2304
rect 9582 2292 9588 2304
rect 9364 2264 9588 2292
rect 9364 2252 9370 2264
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 14274 2292 14280 2304
rect 14235 2264 14280 2292
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 1104 2202 28336 2224
rect 1104 2150 1782 2202
rect 1834 2150 1846 2202
rect 1898 2150 1910 2202
rect 1962 2150 1974 2202
rect 2026 2150 4782 2202
rect 4834 2150 4846 2202
rect 4898 2150 4910 2202
rect 4962 2150 4974 2202
rect 5026 2150 7782 2202
rect 7834 2150 7846 2202
rect 7898 2150 7910 2202
rect 7962 2150 7974 2202
rect 8026 2150 10782 2202
rect 10834 2150 10846 2202
rect 10898 2150 10910 2202
rect 10962 2150 10974 2202
rect 11026 2150 13782 2202
rect 13834 2150 13846 2202
rect 13898 2150 13910 2202
rect 13962 2150 13974 2202
rect 14026 2150 16782 2202
rect 16834 2150 16846 2202
rect 16898 2150 16910 2202
rect 16962 2150 16974 2202
rect 17026 2150 19782 2202
rect 19834 2150 19846 2202
rect 19898 2150 19910 2202
rect 19962 2150 19974 2202
rect 20026 2150 22782 2202
rect 22834 2150 22846 2202
rect 22898 2150 22910 2202
rect 22962 2150 22974 2202
rect 23026 2150 25782 2202
rect 25834 2150 25846 2202
rect 25898 2150 25910 2202
rect 25962 2150 25974 2202
rect 26026 2150 28336 2202
rect 1104 2128 28336 2150
rect 14 8 20 60
rect 72 48 78 60
rect 9950 48 9956 60
rect 72 20 9956 48
rect 72 8 78 20
rect 9950 8 9956 20
rect 10008 8 10014 60
<< via1 >>
rect 1782 29350 1834 29402
rect 1846 29350 1898 29402
rect 1910 29350 1962 29402
rect 1974 29350 2026 29402
rect 4782 29350 4834 29402
rect 4846 29350 4898 29402
rect 4910 29350 4962 29402
rect 4974 29350 5026 29402
rect 7782 29350 7834 29402
rect 7846 29350 7898 29402
rect 7910 29350 7962 29402
rect 7974 29350 8026 29402
rect 10782 29350 10834 29402
rect 10846 29350 10898 29402
rect 10910 29350 10962 29402
rect 10974 29350 11026 29402
rect 13782 29350 13834 29402
rect 13846 29350 13898 29402
rect 13910 29350 13962 29402
rect 13974 29350 14026 29402
rect 16782 29350 16834 29402
rect 16846 29350 16898 29402
rect 16910 29350 16962 29402
rect 16974 29350 17026 29402
rect 19782 29350 19834 29402
rect 19846 29350 19898 29402
rect 19910 29350 19962 29402
rect 19974 29350 20026 29402
rect 22782 29350 22834 29402
rect 22846 29350 22898 29402
rect 22910 29350 22962 29402
rect 22974 29350 23026 29402
rect 25782 29350 25834 29402
rect 25846 29350 25898 29402
rect 25910 29350 25962 29402
rect 25974 29350 26026 29402
rect 3282 28806 3334 28858
rect 3346 28806 3398 28858
rect 3410 28806 3462 28858
rect 3474 28806 3526 28858
rect 6282 28806 6334 28858
rect 6346 28806 6398 28858
rect 6410 28806 6462 28858
rect 6474 28806 6526 28858
rect 9282 28806 9334 28858
rect 9346 28806 9398 28858
rect 9410 28806 9462 28858
rect 9474 28806 9526 28858
rect 12282 28806 12334 28858
rect 12346 28806 12398 28858
rect 12410 28806 12462 28858
rect 12474 28806 12526 28858
rect 15282 28806 15334 28858
rect 15346 28806 15398 28858
rect 15410 28806 15462 28858
rect 15474 28806 15526 28858
rect 18282 28806 18334 28858
rect 18346 28806 18398 28858
rect 18410 28806 18462 28858
rect 18474 28806 18526 28858
rect 21282 28806 21334 28858
rect 21346 28806 21398 28858
rect 21410 28806 21462 28858
rect 21474 28806 21526 28858
rect 24282 28806 24334 28858
rect 24346 28806 24398 28858
rect 24410 28806 24462 28858
rect 24474 28806 24526 28858
rect 27282 28806 27334 28858
rect 27346 28806 27398 28858
rect 27410 28806 27462 28858
rect 27474 28806 27526 28858
rect 1782 28262 1834 28314
rect 1846 28262 1898 28314
rect 1910 28262 1962 28314
rect 1974 28262 2026 28314
rect 4782 28262 4834 28314
rect 4846 28262 4898 28314
rect 4910 28262 4962 28314
rect 4974 28262 5026 28314
rect 7782 28262 7834 28314
rect 7846 28262 7898 28314
rect 7910 28262 7962 28314
rect 7974 28262 8026 28314
rect 10782 28262 10834 28314
rect 10846 28262 10898 28314
rect 10910 28262 10962 28314
rect 10974 28262 11026 28314
rect 13782 28262 13834 28314
rect 13846 28262 13898 28314
rect 13910 28262 13962 28314
rect 13974 28262 14026 28314
rect 16782 28262 16834 28314
rect 16846 28262 16898 28314
rect 16910 28262 16962 28314
rect 16974 28262 17026 28314
rect 19782 28262 19834 28314
rect 19846 28262 19898 28314
rect 19910 28262 19962 28314
rect 19974 28262 20026 28314
rect 22782 28262 22834 28314
rect 22846 28262 22898 28314
rect 22910 28262 22962 28314
rect 22974 28262 23026 28314
rect 25782 28262 25834 28314
rect 25846 28262 25898 28314
rect 25910 28262 25962 28314
rect 25974 28262 26026 28314
rect 3282 27718 3334 27770
rect 3346 27718 3398 27770
rect 3410 27718 3462 27770
rect 3474 27718 3526 27770
rect 6282 27718 6334 27770
rect 6346 27718 6398 27770
rect 6410 27718 6462 27770
rect 6474 27718 6526 27770
rect 9282 27718 9334 27770
rect 9346 27718 9398 27770
rect 9410 27718 9462 27770
rect 9474 27718 9526 27770
rect 12282 27718 12334 27770
rect 12346 27718 12398 27770
rect 12410 27718 12462 27770
rect 12474 27718 12526 27770
rect 15282 27718 15334 27770
rect 15346 27718 15398 27770
rect 15410 27718 15462 27770
rect 15474 27718 15526 27770
rect 18282 27718 18334 27770
rect 18346 27718 18398 27770
rect 18410 27718 18462 27770
rect 18474 27718 18526 27770
rect 21282 27718 21334 27770
rect 21346 27718 21398 27770
rect 21410 27718 21462 27770
rect 21474 27718 21526 27770
rect 24282 27718 24334 27770
rect 24346 27718 24398 27770
rect 24410 27718 24462 27770
rect 24474 27718 24526 27770
rect 27282 27718 27334 27770
rect 27346 27718 27398 27770
rect 27410 27718 27462 27770
rect 27474 27718 27526 27770
rect 23112 27412 23164 27464
rect 24584 27412 24636 27464
rect 21640 27344 21692 27396
rect 1782 27174 1834 27226
rect 1846 27174 1898 27226
rect 1910 27174 1962 27226
rect 1974 27174 2026 27226
rect 4782 27174 4834 27226
rect 4846 27174 4898 27226
rect 4910 27174 4962 27226
rect 4974 27174 5026 27226
rect 7782 27174 7834 27226
rect 7846 27174 7898 27226
rect 7910 27174 7962 27226
rect 7974 27174 8026 27226
rect 10782 27174 10834 27226
rect 10846 27174 10898 27226
rect 10910 27174 10962 27226
rect 10974 27174 11026 27226
rect 13782 27174 13834 27226
rect 13846 27174 13898 27226
rect 13910 27174 13962 27226
rect 13974 27174 14026 27226
rect 16782 27174 16834 27226
rect 16846 27174 16898 27226
rect 16910 27174 16962 27226
rect 16974 27174 17026 27226
rect 19782 27174 19834 27226
rect 19846 27174 19898 27226
rect 19910 27174 19962 27226
rect 19974 27174 20026 27226
rect 22782 27174 22834 27226
rect 22846 27174 22898 27226
rect 22910 27174 22962 27226
rect 22974 27174 23026 27226
rect 25782 27174 25834 27226
rect 25846 27174 25898 27226
rect 25910 27174 25962 27226
rect 25974 27174 26026 27226
rect 23112 27115 23164 27124
rect 23112 27081 23121 27115
rect 23121 27081 23155 27115
rect 23155 27081 23164 27115
rect 23112 27072 23164 27081
rect 3282 26630 3334 26682
rect 3346 26630 3398 26682
rect 3410 26630 3462 26682
rect 3474 26630 3526 26682
rect 6282 26630 6334 26682
rect 6346 26630 6398 26682
rect 6410 26630 6462 26682
rect 6474 26630 6526 26682
rect 9282 26630 9334 26682
rect 9346 26630 9398 26682
rect 9410 26630 9462 26682
rect 9474 26630 9526 26682
rect 12282 26630 12334 26682
rect 12346 26630 12398 26682
rect 12410 26630 12462 26682
rect 12474 26630 12526 26682
rect 15282 26630 15334 26682
rect 15346 26630 15398 26682
rect 15410 26630 15462 26682
rect 15474 26630 15526 26682
rect 18282 26630 18334 26682
rect 18346 26630 18398 26682
rect 18410 26630 18462 26682
rect 18474 26630 18526 26682
rect 21282 26630 21334 26682
rect 21346 26630 21398 26682
rect 21410 26630 21462 26682
rect 21474 26630 21526 26682
rect 24282 26630 24334 26682
rect 24346 26630 24398 26682
rect 24410 26630 24462 26682
rect 24474 26630 24526 26682
rect 27282 26630 27334 26682
rect 27346 26630 27398 26682
rect 27410 26630 27462 26682
rect 27474 26630 27526 26682
rect 1782 26086 1834 26138
rect 1846 26086 1898 26138
rect 1910 26086 1962 26138
rect 1974 26086 2026 26138
rect 4782 26086 4834 26138
rect 4846 26086 4898 26138
rect 4910 26086 4962 26138
rect 4974 26086 5026 26138
rect 7782 26086 7834 26138
rect 7846 26086 7898 26138
rect 7910 26086 7962 26138
rect 7974 26086 8026 26138
rect 10782 26086 10834 26138
rect 10846 26086 10898 26138
rect 10910 26086 10962 26138
rect 10974 26086 11026 26138
rect 13782 26086 13834 26138
rect 13846 26086 13898 26138
rect 13910 26086 13962 26138
rect 13974 26086 14026 26138
rect 16782 26086 16834 26138
rect 16846 26086 16898 26138
rect 16910 26086 16962 26138
rect 16974 26086 17026 26138
rect 19782 26086 19834 26138
rect 19846 26086 19898 26138
rect 19910 26086 19962 26138
rect 19974 26086 20026 26138
rect 22782 26086 22834 26138
rect 22846 26086 22898 26138
rect 22910 26086 22962 26138
rect 22974 26086 23026 26138
rect 25782 26086 25834 26138
rect 25846 26086 25898 26138
rect 25910 26086 25962 26138
rect 25974 26086 26026 26138
rect 3282 25542 3334 25594
rect 3346 25542 3398 25594
rect 3410 25542 3462 25594
rect 3474 25542 3526 25594
rect 6282 25542 6334 25594
rect 6346 25542 6398 25594
rect 6410 25542 6462 25594
rect 6474 25542 6526 25594
rect 9282 25542 9334 25594
rect 9346 25542 9398 25594
rect 9410 25542 9462 25594
rect 9474 25542 9526 25594
rect 12282 25542 12334 25594
rect 12346 25542 12398 25594
rect 12410 25542 12462 25594
rect 12474 25542 12526 25594
rect 15282 25542 15334 25594
rect 15346 25542 15398 25594
rect 15410 25542 15462 25594
rect 15474 25542 15526 25594
rect 18282 25542 18334 25594
rect 18346 25542 18398 25594
rect 18410 25542 18462 25594
rect 18474 25542 18526 25594
rect 21282 25542 21334 25594
rect 21346 25542 21398 25594
rect 21410 25542 21462 25594
rect 21474 25542 21526 25594
rect 24282 25542 24334 25594
rect 24346 25542 24398 25594
rect 24410 25542 24462 25594
rect 24474 25542 24526 25594
rect 27282 25542 27334 25594
rect 27346 25542 27398 25594
rect 27410 25542 27462 25594
rect 27474 25542 27526 25594
rect 1782 24998 1834 25050
rect 1846 24998 1898 25050
rect 1910 24998 1962 25050
rect 1974 24998 2026 25050
rect 4782 24998 4834 25050
rect 4846 24998 4898 25050
rect 4910 24998 4962 25050
rect 4974 24998 5026 25050
rect 7782 24998 7834 25050
rect 7846 24998 7898 25050
rect 7910 24998 7962 25050
rect 7974 24998 8026 25050
rect 10782 24998 10834 25050
rect 10846 24998 10898 25050
rect 10910 24998 10962 25050
rect 10974 24998 11026 25050
rect 13782 24998 13834 25050
rect 13846 24998 13898 25050
rect 13910 24998 13962 25050
rect 13974 24998 14026 25050
rect 16782 24998 16834 25050
rect 16846 24998 16898 25050
rect 16910 24998 16962 25050
rect 16974 24998 17026 25050
rect 19782 24998 19834 25050
rect 19846 24998 19898 25050
rect 19910 24998 19962 25050
rect 19974 24998 20026 25050
rect 22782 24998 22834 25050
rect 22846 24998 22898 25050
rect 22910 24998 22962 25050
rect 22974 24998 23026 25050
rect 25782 24998 25834 25050
rect 25846 24998 25898 25050
rect 25910 24998 25962 25050
rect 25974 24998 26026 25050
rect 3282 24454 3334 24506
rect 3346 24454 3398 24506
rect 3410 24454 3462 24506
rect 3474 24454 3526 24506
rect 6282 24454 6334 24506
rect 6346 24454 6398 24506
rect 6410 24454 6462 24506
rect 6474 24454 6526 24506
rect 9282 24454 9334 24506
rect 9346 24454 9398 24506
rect 9410 24454 9462 24506
rect 9474 24454 9526 24506
rect 12282 24454 12334 24506
rect 12346 24454 12398 24506
rect 12410 24454 12462 24506
rect 12474 24454 12526 24506
rect 15282 24454 15334 24506
rect 15346 24454 15398 24506
rect 15410 24454 15462 24506
rect 15474 24454 15526 24506
rect 18282 24454 18334 24506
rect 18346 24454 18398 24506
rect 18410 24454 18462 24506
rect 18474 24454 18526 24506
rect 21282 24454 21334 24506
rect 21346 24454 21398 24506
rect 21410 24454 21462 24506
rect 21474 24454 21526 24506
rect 24282 24454 24334 24506
rect 24346 24454 24398 24506
rect 24410 24454 24462 24506
rect 24474 24454 24526 24506
rect 27282 24454 27334 24506
rect 27346 24454 27398 24506
rect 27410 24454 27462 24506
rect 27474 24454 27526 24506
rect 1782 23910 1834 23962
rect 1846 23910 1898 23962
rect 1910 23910 1962 23962
rect 1974 23910 2026 23962
rect 4782 23910 4834 23962
rect 4846 23910 4898 23962
rect 4910 23910 4962 23962
rect 4974 23910 5026 23962
rect 7782 23910 7834 23962
rect 7846 23910 7898 23962
rect 7910 23910 7962 23962
rect 7974 23910 8026 23962
rect 10782 23910 10834 23962
rect 10846 23910 10898 23962
rect 10910 23910 10962 23962
rect 10974 23910 11026 23962
rect 13782 23910 13834 23962
rect 13846 23910 13898 23962
rect 13910 23910 13962 23962
rect 13974 23910 14026 23962
rect 16782 23910 16834 23962
rect 16846 23910 16898 23962
rect 16910 23910 16962 23962
rect 16974 23910 17026 23962
rect 19782 23910 19834 23962
rect 19846 23910 19898 23962
rect 19910 23910 19962 23962
rect 19974 23910 20026 23962
rect 22782 23910 22834 23962
rect 22846 23910 22898 23962
rect 22910 23910 22962 23962
rect 22974 23910 23026 23962
rect 25782 23910 25834 23962
rect 25846 23910 25898 23962
rect 25910 23910 25962 23962
rect 25974 23910 26026 23962
rect 3282 23366 3334 23418
rect 3346 23366 3398 23418
rect 3410 23366 3462 23418
rect 3474 23366 3526 23418
rect 6282 23366 6334 23418
rect 6346 23366 6398 23418
rect 6410 23366 6462 23418
rect 6474 23366 6526 23418
rect 9282 23366 9334 23418
rect 9346 23366 9398 23418
rect 9410 23366 9462 23418
rect 9474 23366 9526 23418
rect 12282 23366 12334 23418
rect 12346 23366 12398 23418
rect 12410 23366 12462 23418
rect 12474 23366 12526 23418
rect 15282 23366 15334 23418
rect 15346 23366 15398 23418
rect 15410 23366 15462 23418
rect 15474 23366 15526 23418
rect 18282 23366 18334 23418
rect 18346 23366 18398 23418
rect 18410 23366 18462 23418
rect 18474 23366 18526 23418
rect 21282 23366 21334 23418
rect 21346 23366 21398 23418
rect 21410 23366 21462 23418
rect 21474 23366 21526 23418
rect 24282 23366 24334 23418
rect 24346 23366 24398 23418
rect 24410 23366 24462 23418
rect 24474 23366 24526 23418
rect 27282 23366 27334 23418
rect 27346 23366 27398 23418
rect 27410 23366 27462 23418
rect 27474 23366 27526 23418
rect 1782 22822 1834 22874
rect 1846 22822 1898 22874
rect 1910 22822 1962 22874
rect 1974 22822 2026 22874
rect 4782 22822 4834 22874
rect 4846 22822 4898 22874
rect 4910 22822 4962 22874
rect 4974 22822 5026 22874
rect 7782 22822 7834 22874
rect 7846 22822 7898 22874
rect 7910 22822 7962 22874
rect 7974 22822 8026 22874
rect 10782 22822 10834 22874
rect 10846 22822 10898 22874
rect 10910 22822 10962 22874
rect 10974 22822 11026 22874
rect 13782 22822 13834 22874
rect 13846 22822 13898 22874
rect 13910 22822 13962 22874
rect 13974 22822 14026 22874
rect 16782 22822 16834 22874
rect 16846 22822 16898 22874
rect 16910 22822 16962 22874
rect 16974 22822 17026 22874
rect 19782 22822 19834 22874
rect 19846 22822 19898 22874
rect 19910 22822 19962 22874
rect 19974 22822 20026 22874
rect 22782 22822 22834 22874
rect 22846 22822 22898 22874
rect 22910 22822 22962 22874
rect 22974 22822 23026 22874
rect 25782 22822 25834 22874
rect 25846 22822 25898 22874
rect 25910 22822 25962 22874
rect 25974 22822 26026 22874
rect 3282 22278 3334 22330
rect 3346 22278 3398 22330
rect 3410 22278 3462 22330
rect 3474 22278 3526 22330
rect 6282 22278 6334 22330
rect 6346 22278 6398 22330
rect 6410 22278 6462 22330
rect 6474 22278 6526 22330
rect 9282 22278 9334 22330
rect 9346 22278 9398 22330
rect 9410 22278 9462 22330
rect 9474 22278 9526 22330
rect 12282 22278 12334 22330
rect 12346 22278 12398 22330
rect 12410 22278 12462 22330
rect 12474 22278 12526 22330
rect 15282 22278 15334 22330
rect 15346 22278 15398 22330
rect 15410 22278 15462 22330
rect 15474 22278 15526 22330
rect 18282 22278 18334 22330
rect 18346 22278 18398 22330
rect 18410 22278 18462 22330
rect 18474 22278 18526 22330
rect 21282 22278 21334 22330
rect 21346 22278 21398 22330
rect 21410 22278 21462 22330
rect 21474 22278 21526 22330
rect 24282 22278 24334 22330
rect 24346 22278 24398 22330
rect 24410 22278 24462 22330
rect 24474 22278 24526 22330
rect 27282 22278 27334 22330
rect 27346 22278 27398 22330
rect 27410 22278 27462 22330
rect 27474 22278 27526 22330
rect 1782 21734 1834 21786
rect 1846 21734 1898 21786
rect 1910 21734 1962 21786
rect 1974 21734 2026 21786
rect 4782 21734 4834 21786
rect 4846 21734 4898 21786
rect 4910 21734 4962 21786
rect 4974 21734 5026 21786
rect 7782 21734 7834 21786
rect 7846 21734 7898 21786
rect 7910 21734 7962 21786
rect 7974 21734 8026 21786
rect 10782 21734 10834 21786
rect 10846 21734 10898 21786
rect 10910 21734 10962 21786
rect 10974 21734 11026 21786
rect 13782 21734 13834 21786
rect 13846 21734 13898 21786
rect 13910 21734 13962 21786
rect 13974 21734 14026 21786
rect 16782 21734 16834 21786
rect 16846 21734 16898 21786
rect 16910 21734 16962 21786
rect 16974 21734 17026 21786
rect 19782 21734 19834 21786
rect 19846 21734 19898 21786
rect 19910 21734 19962 21786
rect 19974 21734 20026 21786
rect 22782 21734 22834 21786
rect 22846 21734 22898 21786
rect 22910 21734 22962 21786
rect 22974 21734 23026 21786
rect 25782 21734 25834 21786
rect 25846 21734 25898 21786
rect 25910 21734 25962 21786
rect 25974 21734 26026 21786
rect 3282 21190 3334 21242
rect 3346 21190 3398 21242
rect 3410 21190 3462 21242
rect 3474 21190 3526 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 6410 21190 6462 21242
rect 6474 21190 6526 21242
rect 9282 21190 9334 21242
rect 9346 21190 9398 21242
rect 9410 21190 9462 21242
rect 9474 21190 9526 21242
rect 12282 21190 12334 21242
rect 12346 21190 12398 21242
rect 12410 21190 12462 21242
rect 12474 21190 12526 21242
rect 15282 21190 15334 21242
rect 15346 21190 15398 21242
rect 15410 21190 15462 21242
rect 15474 21190 15526 21242
rect 18282 21190 18334 21242
rect 18346 21190 18398 21242
rect 18410 21190 18462 21242
rect 18474 21190 18526 21242
rect 21282 21190 21334 21242
rect 21346 21190 21398 21242
rect 21410 21190 21462 21242
rect 21474 21190 21526 21242
rect 24282 21190 24334 21242
rect 24346 21190 24398 21242
rect 24410 21190 24462 21242
rect 24474 21190 24526 21242
rect 27282 21190 27334 21242
rect 27346 21190 27398 21242
rect 27410 21190 27462 21242
rect 27474 21190 27526 21242
rect 1782 20646 1834 20698
rect 1846 20646 1898 20698
rect 1910 20646 1962 20698
rect 1974 20646 2026 20698
rect 4782 20646 4834 20698
rect 4846 20646 4898 20698
rect 4910 20646 4962 20698
rect 4974 20646 5026 20698
rect 7782 20646 7834 20698
rect 7846 20646 7898 20698
rect 7910 20646 7962 20698
rect 7974 20646 8026 20698
rect 10782 20646 10834 20698
rect 10846 20646 10898 20698
rect 10910 20646 10962 20698
rect 10974 20646 11026 20698
rect 13782 20646 13834 20698
rect 13846 20646 13898 20698
rect 13910 20646 13962 20698
rect 13974 20646 14026 20698
rect 16782 20646 16834 20698
rect 16846 20646 16898 20698
rect 16910 20646 16962 20698
rect 16974 20646 17026 20698
rect 19782 20646 19834 20698
rect 19846 20646 19898 20698
rect 19910 20646 19962 20698
rect 19974 20646 20026 20698
rect 22782 20646 22834 20698
rect 22846 20646 22898 20698
rect 22910 20646 22962 20698
rect 22974 20646 23026 20698
rect 25782 20646 25834 20698
rect 25846 20646 25898 20698
rect 25910 20646 25962 20698
rect 25974 20646 26026 20698
rect 3282 20102 3334 20154
rect 3346 20102 3398 20154
rect 3410 20102 3462 20154
rect 3474 20102 3526 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 6410 20102 6462 20154
rect 6474 20102 6526 20154
rect 9282 20102 9334 20154
rect 9346 20102 9398 20154
rect 9410 20102 9462 20154
rect 9474 20102 9526 20154
rect 12282 20102 12334 20154
rect 12346 20102 12398 20154
rect 12410 20102 12462 20154
rect 12474 20102 12526 20154
rect 15282 20102 15334 20154
rect 15346 20102 15398 20154
rect 15410 20102 15462 20154
rect 15474 20102 15526 20154
rect 18282 20102 18334 20154
rect 18346 20102 18398 20154
rect 18410 20102 18462 20154
rect 18474 20102 18526 20154
rect 21282 20102 21334 20154
rect 21346 20102 21398 20154
rect 21410 20102 21462 20154
rect 21474 20102 21526 20154
rect 24282 20102 24334 20154
rect 24346 20102 24398 20154
rect 24410 20102 24462 20154
rect 24474 20102 24526 20154
rect 27282 20102 27334 20154
rect 27346 20102 27398 20154
rect 27410 20102 27462 20154
rect 27474 20102 27526 20154
rect 1782 19558 1834 19610
rect 1846 19558 1898 19610
rect 1910 19558 1962 19610
rect 1974 19558 2026 19610
rect 4782 19558 4834 19610
rect 4846 19558 4898 19610
rect 4910 19558 4962 19610
rect 4974 19558 5026 19610
rect 7782 19558 7834 19610
rect 7846 19558 7898 19610
rect 7910 19558 7962 19610
rect 7974 19558 8026 19610
rect 10782 19558 10834 19610
rect 10846 19558 10898 19610
rect 10910 19558 10962 19610
rect 10974 19558 11026 19610
rect 13782 19558 13834 19610
rect 13846 19558 13898 19610
rect 13910 19558 13962 19610
rect 13974 19558 14026 19610
rect 16782 19558 16834 19610
rect 16846 19558 16898 19610
rect 16910 19558 16962 19610
rect 16974 19558 17026 19610
rect 19782 19558 19834 19610
rect 19846 19558 19898 19610
rect 19910 19558 19962 19610
rect 19974 19558 20026 19610
rect 22782 19558 22834 19610
rect 22846 19558 22898 19610
rect 22910 19558 22962 19610
rect 22974 19558 23026 19610
rect 25782 19558 25834 19610
rect 25846 19558 25898 19610
rect 25910 19558 25962 19610
rect 25974 19558 26026 19610
rect 3282 19014 3334 19066
rect 3346 19014 3398 19066
rect 3410 19014 3462 19066
rect 3474 19014 3526 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 6410 19014 6462 19066
rect 6474 19014 6526 19066
rect 9282 19014 9334 19066
rect 9346 19014 9398 19066
rect 9410 19014 9462 19066
rect 9474 19014 9526 19066
rect 12282 19014 12334 19066
rect 12346 19014 12398 19066
rect 12410 19014 12462 19066
rect 12474 19014 12526 19066
rect 15282 19014 15334 19066
rect 15346 19014 15398 19066
rect 15410 19014 15462 19066
rect 15474 19014 15526 19066
rect 18282 19014 18334 19066
rect 18346 19014 18398 19066
rect 18410 19014 18462 19066
rect 18474 19014 18526 19066
rect 21282 19014 21334 19066
rect 21346 19014 21398 19066
rect 21410 19014 21462 19066
rect 21474 19014 21526 19066
rect 24282 19014 24334 19066
rect 24346 19014 24398 19066
rect 24410 19014 24462 19066
rect 24474 19014 24526 19066
rect 27282 19014 27334 19066
rect 27346 19014 27398 19066
rect 27410 19014 27462 19066
rect 27474 19014 27526 19066
rect 1782 18470 1834 18522
rect 1846 18470 1898 18522
rect 1910 18470 1962 18522
rect 1974 18470 2026 18522
rect 4782 18470 4834 18522
rect 4846 18470 4898 18522
rect 4910 18470 4962 18522
rect 4974 18470 5026 18522
rect 7782 18470 7834 18522
rect 7846 18470 7898 18522
rect 7910 18470 7962 18522
rect 7974 18470 8026 18522
rect 10782 18470 10834 18522
rect 10846 18470 10898 18522
rect 10910 18470 10962 18522
rect 10974 18470 11026 18522
rect 13782 18470 13834 18522
rect 13846 18470 13898 18522
rect 13910 18470 13962 18522
rect 13974 18470 14026 18522
rect 16782 18470 16834 18522
rect 16846 18470 16898 18522
rect 16910 18470 16962 18522
rect 16974 18470 17026 18522
rect 19782 18470 19834 18522
rect 19846 18470 19898 18522
rect 19910 18470 19962 18522
rect 19974 18470 20026 18522
rect 22782 18470 22834 18522
rect 22846 18470 22898 18522
rect 22910 18470 22962 18522
rect 22974 18470 23026 18522
rect 25782 18470 25834 18522
rect 25846 18470 25898 18522
rect 25910 18470 25962 18522
rect 25974 18470 26026 18522
rect 3282 17926 3334 17978
rect 3346 17926 3398 17978
rect 3410 17926 3462 17978
rect 3474 17926 3526 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 6410 17926 6462 17978
rect 6474 17926 6526 17978
rect 9282 17926 9334 17978
rect 9346 17926 9398 17978
rect 9410 17926 9462 17978
rect 9474 17926 9526 17978
rect 12282 17926 12334 17978
rect 12346 17926 12398 17978
rect 12410 17926 12462 17978
rect 12474 17926 12526 17978
rect 15282 17926 15334 17978
rect 15346 17926 15398 17978
rect 15410 17926 15462 17978
rect 15474 17926 15526 17978
rect 18282 17926 18334 17978
rect 18346 17926 18398 17978
rect 18410 17926 18462 17978
rect 18474 17926 18526 17978
rect 21282 17926 21334 17978
rect 21346 17926 21398 17978
rect 21410 17926 21462 17978
rect 21474 17926 21526 17978
rect 24282 17926 24334 17978
rect 24346 17926 24398 17978
rect 24410 17926 24462 17978
rect 24474 17926 24526 17978
rect 27282 17926 27334 17978
rect 27346 17926 27398 17978
rect 27410 17926 27462 17978
rect 27474 17926 27526 17978
rect 1782 17382 1834 17434
rect 1846 17382 1898 17434
rect 1910 17382 1962 17434
rect 1974 17382 2026 17434
rect 4782 17382 4834 17434
rect 4846 17382 4898 17434
rect 4910 17382 4962 17434
rect 4974 17382 5026 17434
rect 7782 17382 7834 17434
rect 7846 17382 7898 17434
rect 7910 17382 7962 17434
rect 7974 17382 8026 17434
rect 10782 17382 10834 17434
rect 10846 17382 10898 17434
rect 10910 17382 10962 17434
rect 10974 17382 11026 17434
rect 13782 17382 13834 17434
rect 13846 17382 13898 17434
rect 13910 17382 13962 17434
rect 13974 17382 14026 17434
rect 16782 17382 16834 17434
rect 16846 17382 16898 17434
rect 16910 17382 16962 17434
rect 16974 17382 17026 17434
rect 19782 17382 19834 17434
rect 19846 17382 19898 17434
rect 19910 17382 19962 17434
rect 19974 17382 20026 17434
rect 22782 17382 22834 17434
rect 22846 17382 22898 17434
rect 22910 17382 22962 17434
rect 22974 17382 23026 17434
rect 25782 17382 25834 17434
rect 25846 17382 25898 17434
rect 25910 17382 25962 17434
rect 25974 17382 26026 17434
rect 3282 16838 3334 16890
rect 3346 16838 3398 16890
rect 3410 16838 3462 16890
rect 3474 16838 3526 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 6410 16838 6462 16890
rect 6474 16838 6526 16890
rect 9282 16838 9334 16890
rect 9346 16838 9398 16890
rect 9410 16838 9462 16890
rect 9474 16838 9526 16890
rect 12282 16838 12334 16890
rect 12346 16838 12398 16890
rect 12410 16838 12462 16890
rect 12474 16838 12526 16890
rect 15282 16838 15334 16890
rect 15346 16838 15398 16890
rect 15410 16838 15462 16890
rect 15474 16838 15526 16890
rect 18282 16838 18334 16890
rect 18346 16838 18398 16890
rect 18410 16838 18462 16890
rect 18474 16838 18526 16890
rect 21282 16838 21334 16890
rect 21346 16838 21398 16890
rect 21410 16838 21462 16890
rect 21474 16838 21526 16890
rect 24282 16838 24334 16890
rect 24346 16838 24398 16890
rect 24410 16838 24462 16890
rect 24474 16838 24526 16890
rect 27282 16838 27334 16890
rect 27346 16838 27398 16890
rect 27410 16838 27462 16890
rect 27474 16838 27526 16890
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 15568 16532 15620 16584
rect 15752 16464 15804 16516
rect 16488 16464 16540 16516
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 14924 16396 14976 16448
rect 1782 16294 1834 16346
rect 1846 16294 1898 16346
rect 1910 16294 1962 16346
rect 1974 16294 2026 16346
rect 4782 16294 4834 16346
rect 4846 16294 4898 16346
rect 4910 16294 4962 16346
rect 4974 16294 5026 16346
rect 7782 16294 7834 16346
rect 7846 16294 7898 16346
rect 7910 16294 7962 16346
rect 7974 16294 8026 16346
rect 10782 16294 10834 16346
rect 10846 16294 10898 16346
rect 10910 16294 10962 16346
rect 10974 16294 11026 16346
rect 13782 16294 13834 16346
rect 13846 16294 13898 16346
rect 13910 16294 13962 16346
rect 13974 16294 14026 16346
rect 16782 16294 16834 16346
rect 16846 16294 16898 16346
rect 16910 16294 16962 16346
rect 16974 16294 17026 16346
rect 19782 16294 19834 16346
rect 19846 16294 19898 16346
rect 19910 16294 19962 16346
rect 19974 16294 20026 16346
rect 22782 16294 22834 16346
rect 22846 16294 22898 16346
rect 22910 16294 22962 16346
rect 22974 16294 23026 16346
rect 25782 16294 25834 16346
rect 25846 16294 25898 16346
rect 25910 16294 25962 16346
rect 25974 16294 26026 16346
rect 14924 16124 14976 16176
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 14556 15988 14608 16040
rect 15660 15988 15712 16040
rect 15568 15920 15620 15972
rect 14096 15852 14148 15904
rect 16580 15852 16632 15904
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 3282 15750 3334 15802
rect 3346 15750 3398 15802
rect 3410 15750 3462 15802
rect 3474 15750 3526 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 6410 15750 6462 15802
rect 6474 15750 6526 15802
rect 9282 15750 9334 15802
rect 9346 15750 9398 15802
rect 9410 15750 9462 15802
rect 9474 15750 9526 15802
rect 12282 15750 12334 15802
rect 12346 15750 12398 15802
rect 12410 15750 12462 15802
rect 12474 15750 12526 15802
rect 15282 15750 15334 15802
rect 15346 15750 15398 15802
rect 15410 15750 15462 15802
rect 15474 15750 15526 15802
rect 18282 15750 18334 15802
rect 18346 15750 18398 15802
rect 18410 15750 18462 15802
rect 18474 15750 18526 15802
rect 21282 15750 21334 15802
rect 21346 15750 21398 15802
rect 21410 15750 21462 15802
rect 21474 15750 21526 15802
rect 24282 15750 24334 15802
rect 24346 15750 24398 15802
rect 24410 15750 24462 15802
rect 24474 15750 24526 15802
rect 27282 15750 27334 15802
rect 27346 15750 27398 15802
rect 27410 15750 27462 15802
rect 27474 15750 27526 15802
rect 14280 15648 14332 15700
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 15384 15444 15436 15496
rect 15752 15580 15804 15632
rect 16580 15580 16632 15632
rect 16212 15512 16264 15564
rect 15476 15419 15528 15428
rect 15476 15385 15485 15419
rect 15485 15385 15519 15419
rect 15519 15385 15528 15419
rect 15476 15376 15528 15385
rect 16028 15419 16080 15428
rect 16028 15385 16037 15419
rect 16037 15385 16071 15419
rect 16071 15385 16080 15419
rect 16028 15376 16080 15385
rect 17316 15444 17368 15496
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 18144 15444 18196 15496
rect 18512 15444 18564 15496
rect 20536 15444 20588 15496
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 16396 15351 16448 15360
rect 16396 15317 16405 15351
rect 16405 15317 16439 15351
rect 16439 15317 16448 15351
rect 16396 15308 16448 15317
rect 18788 15308 18840 15360
rect 19156 15308 19208 15360
rect 1782 15206 1834 15258
rect 1846 15206 1898 15258
rect 1910 15206 1962 15258
rect 1974 15206 2026 15258
rect 4782 15206 4834 15258
rect 4846 15206 4898 15258
rect 4910 15206 4962 15258
rect 4974 15206 5026 15258
rect 7782 15206 7834 15258
rect 7846 15206 7898 15258
rect 7910 15206 7962 15258
rect 7974 15206 8026 15258
rect 10782 15206 10834 15258
rect 10846 15206 10898 15258
rect 10910 15206 10962 15258
rect 10974 15206 11026 15258
rect 13782 15206 13834 15258
rect 13846 15206 13898 15258
rect 13910 15206 13962 15258
rect 13974 15206 14026 15258
rect 16782 15206 16834 15258
rect 16846 15206 16898 15258
rect 16910 15206 16962 15258
rect 16974 15206 17026 15258
rect 19782 15206 19834 15258
rect 19846 15206 19898 15258
rect 19910 15206 19962 15258
rect 19974 15206 20026 15258
rect 22782 15206 22834 15258
rect 22846 15206 22898 15258
rect 22910 15206 22962 15258
rect 22974 15206 23026 15258
rect 25782 15206 25834 15258
rect 25846 15206 25898 15258
rect 25910 15206 25962 15258
rect 25974 15206 26026 15258
rect 12716 15104 12768 15156
rect 14096 15104 14148 15156
rect 15384 15147 15436 15156
rect 13268 14968 13320 15020
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 17776 15104 17828 15156
rect 14832 15036 14884 15088
rect 15476 15036 15528 15088
rect 14556 14968 14608 15020
rect 15016 14968 15068 15020
rect 15660 14968 15712 15020
rect 16580 15011 16632 15020
rect 16580 14977 16589 15011
rect 16589 14977 16623 15011
rect 16623 14977 16632 15011
rect 16580 14968 16632 14977
rect 17316 15036 17368 15088
rect 17500 15036 17552 15088
rect 18512 15079 18564 15088
rect 18512 15045 18521 15079
rect 18521 15045 18555 15079
rect 18555 15045 18564 15079
rect 18512 15036 18564 15045
rect 18880 15104 18932 15156
rect 21180 15036 21232 15088
rect 18788 14900 18840 14952
rect 19432 14832 19484 14884
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 18144 14764 18196 14816
rect 20352 14943 20404 14952
rect 20352 14909 20361 14943
rect 20361 14909 20395 14943
rect 20395 14909 20404 14943
rect 20352 14900 20404 14909
rect 20628 14943 20680 14952
rect 20628 14909 20637 14943
rect 20637 14909 20671 14943
rect 20671 14909 20680 14943
rect 20628 14900 20680 14909
rect 20720 14764 20772 14816
rect 3282 14662 3334 14714
rect 3346 14662 3398 14714
rect 3410 14662 3462 14714
rect 3474 14662 3526 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 6410 14662 6462 14714
rect 6474 14662 6526 14714
rect 9282 14662 9334 14714
rect 9346 14662 9398 14714
rect 9410 14662 9462 14714
rect 9474 14662 9526 14714
rect 12282 14662 12334 14714
rect 12346 14662 12398 14714
rect 12410 14662 12462 14714
rect 12474 14662 12526 14714
rect 15282 14662 15334 14714
rect 15346 14662 15398 14714
rect 15410 14662 15462 14714
rect 15474 14662 15526 14714
rect 18282 14662 18334 14714
rect 18346 14662 18398 14714
rect 18410 14662 18462 14714
rect 18474 14662 18526 14714
rect 21282 14662 21334 14714
rect 21346 14662 21398 14714
rect 21410 14662 21462 14714
rect 21474 14662 21526 14714
rect 24282 14662 24334 14714
rect 24346 14662 24398 14714
rect 24410 14662 24462 14714
rect 24474 14662 24526 14714
rect 27282 14662 27334 14714
rect 27346 14662 27398 14714
rect 27410 14662 27462 14714
rect 27474 14662 27526 14714
rect 14556 14603 14608 14612
rect 14556 14569 14565 14603
rect 14565 14569 14599 14603
rect 14599 14569 14608 14603
rect 14556 14560 14608 14569
rect 15108 14560 15160 14612
rect 16580 14560 16632 14612
rect 21180 14560 21232 14612
rect 14648 14492 14700 14544
rect 17500 14492 17552 14544
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 14188 14424 14240 14476
rect 15936 14356 15988 14408
rect 16212 14399 16264 14408
rect 16212 14365 16221 14399
rect 16221 14365 16255 14399
rect 16255 14365 16264 14399
rect 16212 14356 16264 14365
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 17132 14356 17184 14408
rect 18788 14399 18840 14408
rect 18788 14365 18797 14399
rect 18797 14365 18831 14399
rect 18831 14365 18840 14399
rect 18788 14356 18840 14365
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 12164 14331 12216 14340
rect 12164 14297 12173 14331
rect 12173 14297 12207 14331
rect 12207 14297 12216 14331
rect 12164 14288 12216 14297
rect 12900 14288 12952 14340
rect 13820 14288 13872 14340
rect 14280 14288 14332 14340
rect 19432 14356 19484 14408
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 20628 14288 20680 14340
rect 17960 14263 18012 14272
rect 17960 14229 17969 14263
rect 17969 14229 18003 14263
rect 18003 14229 18012 14263
rect 17960 14220 18012 14229
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 1782 14118 1834 14170
rect 1846 14118 1898 14170
rect 1910 14118 1962 14170
rect 1974 14118 2026 14170
rect 4782 14118 4834 14170
rect 4846 14118 4898 14170
rect 4910 14118 4962 14170
rect 4974 14118 5026 14170
rect 7782 14118 7834 14170
rect 7846 14118 7898 14170
rect 7910 14118 7962 14170
rect 7974 14118 8026 14170
rect 10782 14118 10834 14170
rect 10846 14118 10898 14170
rect 10910 14118 10962 14170
rect 10974 14118 11026 14170
rect 13782 14118 13834 14170
rect 13846 14118 13898 14170
rect 13910 14118 13962 14170
rect 13974 14118 14026 14170
rect 16782 14118 16834 14170
rect 16846 14118 16898 14170
rect 16910 14118 16962 14170
rect 16974 14118 17026 14170
rect 19782 14118 19834 14170
rect 19846 14118 19898 14170
rect 19910 14118 19962 14170
rect 19974 14118 20026 14170
rect 22782 14118 22834 14170
rect 22846 14118 22898 14170
rect 22910 14118 22962 14170
rect 22974 14118 23026 14170
rect 25782 14118 25834 14170
rect 25846 14118 25898 14170
rect 25910 14118 25962 14170
rect 25974 14118 26026 14170
rect 12164 14016 12216 14068
rect 11888 13991 11940 14000
rect 11888 13957 11897 13991
rect 11897 13957 11931 13991
rect 11931 13957 11940 13991
rect 11888 13948 11940 13957
rect 16212 14016 16264 14068
rect 19156 14016 19208 14068
rect 19248 14016 19300 14068
rect 20628 14016 20680 14068
rect 15016 13948 15068 14000
rect 16396 13991 16448 14000
rect 16396 13957 16405 13991
rect 16405 13957 16439 13991
rect 16439 13957 16448 13991
rect 16396 13948 16448 13957
rect 17040 13948 17092 14000
rect 17960 13948 18012 14000
rect 8668 13880 8720 13932
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13452 13923 13504 13932
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 14740 13880 14792 13932
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 15108 13923 15160 13932
rect 14832 13880 14884 13889
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 19064 13923 19116 13932
rect 19064 13889 19073 13923
rect 19073 13889 19107 13923
rect 19107 13889 19116 13923
rect 19064 13880 19116 13889
rect 19156 13880 19208 13932
rect 19524 13880 19576 13932
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 14280 13812 14332 13864
rect 15844 13812 15896 13864
rect 18144 13812 18196 13864
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 12716 13744 12768 13796
rect 13452 13744 13504 13796
rect 13728 13744 13780 13796
rect 16580 13744 16632 13796
rect 20536 13744 20588 13796
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 15752 13676 15804 13728
rect 15936 13676 15988 13728
rect 17132 13676 17184 13728
rect 21180 13676 21232 13728
rect 21640 13676 21692 13728
rect 3282 13574 3334 13626
rect 3346 13574 3398 13626
rect 3410 13574 3462 13626
rect 3474 13574 3526 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 6410 13574 6462 13626
rect 6474 13574 6526 13626
rect 9282 13574 9334 13626
rect 9346 13574 9398 13626
rect 9410 13574 9462 13626
rect 9474 13574 9526 13626
rect 12282 13574 12334 13626
rect 12346 13574 12398 13626
rect 12410 13574 12462 13626
rect 12474 13574 12526 13626
rect 15282 13574 15334 13626
rect 15346 13574 15398 13626
rect 15410 13574 15462 13626
rect 15474 13574 15526 13626
rect 18282 13574 18334 13626
rect 18346 13574 18398 13626
rect 18410 13574 18462 13626
rect 18474 13574 18526 13626
rect 21282 13574 21334 13626
rect 21346 13574 21398 13626
rect 21410 13574 21462 13626
rect 21474 13574 21526 13626
rect 24282 13574 24334 13626
rect 24346 13574 24398 13626
rect 24410 13574 24462 13626
rect 24474 13574 24526 13626
rect 27282 13574 27334 13626
rect 27346 13574 27398 13626
rect 27410 13574 27462 13626
rect 27474 13574 27526 13626
rect 12900 13472 12952 13524
rect 14832 13515 14884 13524
rect 14832 13481 14841 13515
rect 14841 13481 14875 13515
rect 14875 13481 14884 13515
rect 14832 13472 14884 13481
rect 15016 13472 15068 13524
rect 13268 13404 13320 13456
rect 15108 13404 15160 13456
rect 15936 13472 15988 13524
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 13084 13336 13136 13388
rect 14188 13336 14240 13388
rect 14924 13336 14976 13388
rect 13452 13268 13504 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 14280 13268 14332 13320
rect 20904 13404 20956 13456
rect 16672 13336 16724 13388
rect 19340 13336 19392 13388
rect 17040 13311 17092 13320
rect 14740 13200 14792 13252
rect 15660 13200 15712 13252
rect 16212 13243 16264 13252
rect 16212 13209 16221 13243
rect 16221 13209 16255 13243
rect 16255 13209 16264 13243
rect 16212 13200 16264 13209
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 19064 13311 19116 13320
rect 8392 13132 8444 13184
rect 8668 13132 8720 13184
rect 12716 13132 12768 13184
rect 18052 13132 18104 13184
rect 18144 13132 18196 13184
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19156 13268 19208 13320
rect 18880 13200 18932 13252
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 20352 13268 20404 13320
rect 22284 13311 22336 13320
rect 22284 13277 22293 13311
rect 22293 13277 22327 13311
rect 22327 13277 22336 13311
rect 22284 13268 22336 13277
rect 22560 13243 22612 13252
rect 22560 13209 22569 13243
rect 22569 13209 22603 13243
rect 22603 13209 22612 13243
rect 22560 13200 22612 13209
rect 23112 13200 23164 13252
rect 23940 13200 23992 13252
rect 22468 13132 22520 13184
rect 1782 13030 1834 13082
rect 1846 13030 1898 13082
rect 1910 13030 1962 13082
rect 1974 13030 2026 13082
rect 4782 13030 4834 13082
rect 4846 13030 4898 13082
rect 4910 13030 4962 13082
rect 4974 13030 5026 13082
rect 7782 13030 7834 13082
rect 7846 13030 7898 13082
rect 7910 13030 7962 13082
rect 7974 13030 8026 13082
rect 10782 13030 10834 13082
rect 10846 13030 10898 13082
rect 10910 13030 10962 13082
rect 10974 13030 11026 13082
rect 13782 13030 13834 13082
rect 13846 13030 13898 13082
rect 13910 13030 13962 13082
rect 13974 13030 14026 13082
rect 16782 13030 16834 13082
rect 16846 13030 16898 13082
rect 16910 13030 16962 13082
rect 16974 13030 17026 13082
rect 19782 13030 19834 13082
rect 19846 13030 19898 13082
rect 19910 13030 19962 13082
rect 19974 13030 20026 13082
rect 22782 13030 22834 13082
rect 22846 13030 22898 13082
rect 22910 13030 22962 13082
rect 22974 13030 23026 13082
rect 25782 13030 25834 13082
rect 25846 13030 25898 13082
rect 25910 13030 25962 13082
rect 25974 13030 26026 13082
rect 11244 12971 11296 12980
rect 11244 12937 11253 12971
rect 11253 12937 11287 12971
rect 11287 12937 11296 12971
rect 11244 12928 11296 12937
rect 13636 12928 13688 12980
rect 16488 12928 16540 12980
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 14188 12903 14240 12912
rect 14188 12869 14197 12903
rect 14197 12869 14231 12903
rect 14231 12869 14240 12903
rect 17132 12928 17184 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 21732 12928 21784 12980
rect 23112 12928 23164 12980
rect 23940 12971 23992 12980
rect 23940 12937 23949 12971
rect 23949 12937 23983 12971
rect 23983 12937 23992 12971
rect 23940 12928 23992 12937
rect 20168 12903 20220 12912
rect 14188 12860 14240 12869
rect 20168 12869 20177 12903
rect 20177 12869 20211 12903
rect 20211 12869 20220 12903
rect 20168 12860 20220 12869
rect 22284 12860 22336 12912
rect 13268 12835 13320 12844
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 15016 12792 15068 12844
rect 15844 12835 15896 12844
rect 13452 12724 13504 12776
rect 14096 12724 14148 12776
rect 14648 12724 14700 12776
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 19340 12792 19392 12844
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 22468 12792 22520 12844
rect 16488 12724 16540 12776
rect 19156 12724 19208 12776
rect 22652 12767 22704 12776
rect 22652 12733 22661 12767
rect 22661 12733 22695 12767
rect 22695 12733 22704 12767
rect 22652 12724 22704 12733
rect 13544 12656 13596 12708
rect 15568 12656 15620 12708
rect 18696 12656 18748 12708
rect 19616 12656 19668 12708
rect 22560 12656 22612 12708
rect 15108 12588 15160 12640
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 18052 12588 18104 12640
rect 20720 12588 20772 12640
rect 20996 12588 21048 12640
rect 3282 12486 3334 12538
rect 3346 12486 3398 12538
rect 3410 12486 3462 12538
rect 3474 12486 3526 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 6410 12486 6462 12538
rect 6474 12486 6526 12538
rect 9282 12486 9334 12538
rect 9346 12486 9398 12538
rect 9410 12486 9462 12538
rect 9474 12486 9526 12538
rect 12282 12486 12334 12538
rect 12346 12486 12398 12538
rect 12410 12486 12462 12538
rect 12474 12486 12526 12538
rect 15282 12486 15334 12538
rect 15346 12486 15398 12538
rect 15410 12486 15462 12538
rect 15474 12486 15526 12538
rect 18282 12486 18334 12538
rect 18346 12486 18398 12538
rect 18410 12486 18462 12538
rect 18474 12486 18526 12538
rect 21282 12486 21334 12538
rect 21346 12486 21398 12538
rect 21410 12486 21462 12538
rect 21474 12486 21526 12538
rect 24282 12486 24334 12538
rect 24346 12486 24398 12538
rect 24410 12486 24462 12538
rect 24474 12486 24526 12538
rect 27282 12486 27334 12538
rect 27346 12486 27398 12538
rect 27410 12486 27462 12538
rect 27474 12486 27526 12538
rect 8392 12384 8444 12436
rect 13544 12384 13596 12436
rect 15844 12384 15896 12436
rect 20168 12427 20220 12436
rect 15016 12316 15068 12368
rect 16672 12316 16724 12368
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 22560 12427 22612 12436
rect 22560 12393 22569 12427
rect 22569 12393 22603 12427
rect 22603 12393 22612 12427
rect 22560 12384 22612 12393
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 11888 12248 11940 12300
rect 13176 12248 13228 12300
rect 22192 12291 22244 12300
rect 22192 12257 22201 12291
rect 22201 12257 22235 12291
rect 22235 12257 22244 12291
rect 22192 12248 22244 12257
rect 23940 12291 23992 12300
rect 23940 12257 23949 12291
rect 23949 12257 23983 12291
rect 23983 12257 23992 12291
rect 23940 12248 23992 12257
rect 13268 12180 13320 12232
rect 14464 12180 14516 12232
rect 15936 12180 15988 12232
rect 11336 12155 11388 12164
rect 11336 12121 11345 12155
rect 11345 12121 11379 12155
rect 11379 12121 11388 12155
rect 11336 12112 11388 12121
rect 11796 12112 11848 12164
rect 13544 12112 13596 12164
rect 14280 12112 14332 12164
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 17592 12223 17644 12232
rect 16488 12180 16540 12189
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 18144 12180 18196 12232
rect 19156 12180 19208 12232
rect 19524 12180 19576 12232
rect 21732 12223 21784 12232
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 22560 12112 22612 12164
rect 10600 12044 10652 12096
rect 13452 12044 13504 12096
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 14648 12044 14700 12053
rect 18788 12044 18840 12096
rect 19064 12044 19116 12096
rect 21088 12087 21140 12096
rect 21088 12053 21097 12087
rect 21097 12053 21131 12087
rect 21131 12053 21140 12087
rect 21088 12044 21140 12053
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 24308 12044 24360 12096
rect 1782 11942 1834 11994
rect 1846 11942 1898 11994
rect 1910 11942 1962 11994
rect 1974 11942 2026 11994
rect 4782 11942 4834 11994
rect 4846 11942 4898 11994
rect 4910 11942 4962 11994
rect 4974 11942 5026 11994
rect 7782 11942 7834 11994
rect 7846 11942 7898 11994
rect 7910 11942 7962 11994
rect 7974 11942 8026 11994
rect 10782 11942 10834 11994
rect 10846 11942 10898 11994
rect 10910 11942 10962 11994
rect 10974 11942 11026 11994
rect 13782 11942 13834 11994
rect 13846 11942 13898 11994
rect 13910 11942 13962 11994
rect 13974 11942 14026 11994
rect 16782 11942 16834 11994
rect 16846 11942 16898 11994
rect 16910 11942 16962 11994
rect 16974 11942 17026 11994
rect 19782 11942 19834 11994
rect 19846 11942 19898 11994
rect 19910 11942 19962 11994
rect 19974 11942 20026 11994
rect 22782 11942 22834 11994
rect 22846 11942 22898 11994
rect 22910 11942 22962 11994
rect 22974 11942 23026 11994
rect 24308 11951 24360 11960
rect 24308 11917 24317 11951
rect 24317 11917 24351 11951
rect 24351 11917 24360 11951
rect 25782 11942 25834 11994
rect 25846 11942 25898 11994
rect 25910 11942 25962 11994
rect 25974 11942 26026 11994
rect 24308 11908 24360 11917
rect 10600 11840 10652 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 11336 11840 11388 11892
rect 14464 11883 14516 11892
rect 10416 11772 10468 11824
rect 11796 11815 11848 11824
rect 11796 11781 11805 11815
rect 11805 11781 11839 11815
rect 11839 11781 11848 11815
rect 11796 11772 11848 11781
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 16028 11840 16080 11892
rect 8944 11704 8996 11756
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 14188 11772 14240 11824
rect 13452 11747 13504 11756
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 11244 11636 11296 11688
rect 12624 11636 12676 11688
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 15108 11704 15160 11756
rect 15660 11772 15712 11824
rect 17224 11772 17276 11824
rect 17592 11840 17644 11892
rect 22560 11883 22612 11892
rect 17776 11772 17828 11824
rect 22560 11849 22569 11883
rect 22569 11849 22603 11883
rect 22603 11849 22612 11883
rect 22560 11840 22612 11849
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 18696 11747 18748 11756
rect 15568 11704 15620 11713
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 13544 11636 13596 11688
rect 14280 11636 14332 11688
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 13728 11568 13780 11620
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 16488 11636 16540 11688
rect 17132 11636 17184 11688
rect 18052 11636 18104 11688
rect 18420 11679 18472 11688
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 6184 11500 6236 11552
rect 14924 11500 14976 11552
rect 17500 11543 17552 11552
rect 17500 11509 17509 11543
rect 17509 11509 17543 11543
rect 17543 11509 17552 11543
rect 17500 11500 17552 11509
rect 18144 11500 18196 11552
rect 19248 11704 19300 11756
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 21732 11747 21784 11756
rect 19432 11704 19484 11713
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 21732 11713 21741 11747
rect 21741 11713 21775 11747
rect 21775 11713 21784 11747
rect 21732 11704 21784 11713
rect 22284 11704 22336 11756
rect 21824 11636 21876 11688
rect 19800 11611 19852 11620
rect 19800 11577 19809 11611
rect 19809 11577 19843 11611
rect 19843 11577 19852 11611
rect 19800 11568 19852 11577
rect 20996 11568 21048 11620
rect 20352 11543 20404 11552
rect 20352 11509 20361 11543
rect 20361 11509 20395 11543
rect 20395 11509 20404 11543
rect 28724 11636 28776 11688
rect 22284 11543 22336 11552
rect 20352 11500 20404 11509
rect 22284 11509 22293 11543
rect 22293 11509 22327 11543
rect 22327 11509 22336 11543
rect 22284 11500 22336 11509
rect 3282 11398 3334 11450
rect 3346 11398 3398 11450
rect 3410 11398 3462 11450
rect 3474 11398 3526 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 6410 11398 6462 11450
rect 6474 11398 6526 11450
rect 9282 11398 9334 11450
rect 9346 11398 9398 11450
rect 9410 11398 9462 11450
rect 9474 11398 9526 11450
rect 12282 11398 12334 11450
rect 12346 11398 12398 11450
rect 12410 11398 12462 11450
rect 12474 11398 12526 11450
rect 15282 11398 15334 11450
rect 15346 11398 15398 11450
rect 15410 11398 15462 11450
rect 15474 11398 15526 11450
rect 18282 11398 18334 11450
rect 18346 11398 18398 11450
rect 18410 11398 18462 11450
rect 18474 11398 18526 11450
rect 21282 11398 21334 11450
rect 21346 11398 21398 11450
rect 21410 11398 21462 11450
rect 21474 11398 21526 11450
rect 24282 11398 24334 11450
rect 24346 11398 24398 11450
rect 24410 11398 24462 11450
rect 24474 11398 24526 11450
rect 27282 11398 27334 11450
rect 27346 11398 27398 11450
rect 27410 11398 27462 11450
rect 27474 11398 27526 11450
rect 11796 11296 11848 11348
rect 13176 11296 13228 11348
rect 14096 11296 14148 11348
rect 15108 11296 15160 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19248 11296 19300 11348
rect 19524 11339 19576 11348
rect 19524 11305 19533 11339
rect 19533 11305 19567 11339
rect 19567 11305 19576 11339
rect 19524 11296 19576 11305
rect 19800 11296 19852 11348
rect 21088 11296 21140 11348
rect 13728 11271 13780 11280
rect 13728 11237 13737 11271
rect 13737 11237 13771 11271
rect 13771 11237 13780 11271
rect 13728 11228 13780 11237
rect 15660 11228 15712 11280
rect 17224 11228 17276 11280
rect 18788 11271 18840 11280
rect 18788 11237 18797 11271
rect 18797 11237 18831 11271
rect 18831 11237 18840 11271
rect 18788 11228 18840 11237
rect 11336 11160 11388 11212
rect 12716 11160 12768 11212
rect 13452 11160 13504 11212
rect 15016 11160 15068 11212
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8024 11024 8076 11076
rect 9036 11092 9088 11144
rect 11152 11092 11204 11144
rect 11980 11092 12032 11144
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 17592 11160 17644 11212
rect 19616 11203 19668 11212
rect 19616 11169 19625 11203
rect 19625 11169 19659 11203
rect 19659 11169 19668 11203
rect 19616 11160 19668 11169
rect 21824 11203 21876 11212
rect 21824 11169 21833 11203
rect 21833 11169 21867 11203
rect 21867 11169 21876 11203
rect 21824 11160 21876 11169
rect 22284 11160 22336 11212
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 17684 11092 17736 11144
rect 20904 11092 20956 11144
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 15568 11024 15620 11076
rect 16212 11024 16264 11076
rect 21180 11024 21232 11076
rect 22468 11024 22520 11076
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 8944 10956 8996 11008
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 19156 10956 19208 11008
rect 20352 10956 20404 11008
rect 1782 10854 1834 10906
rect 1846 10854 1898 10906
rect 1910 10854 1962 10906
rect 1974 10854 2026 10906
rect 4782 10854 4834 10906
rect 4846 10854 4898 10906
rect 4910 10854 4962 10906
rect 4974 10854 5026 10906
rect 7782 10854 7834 10906
rect 7846 10854 7898 10906
rect 7910 10854 7962 10906
rect 7974 10854 8026 10906
rect 10782 10854 10834 10906
rect 10846 10854 10898 10906
rect 10910 10854 10962 10906
rect 10974 10854 11026 10906
rect 13782 10854 13834 10906
rect 13846 10854 13898 10906
rect 13910 10854 13962 10906
rect 13974 10854 14026 10906
rect 16782 10854 16834 10906
rect 16846 10854 16898 10906
rect 16910 10854 16962 10906
rect 16974 10854 17026 10906
rect 19782 10854 19834 10906
rect 19846 10854 19898 10906
rect 19910 10854 19962 10906
rect 19974 10854 20026 10906
rect 22782 10854 22834 10906
rect 22846 10854 22898 10906
rect 22910 10854 22962 10906
rect 22974 10854 23026 10906
rect 25782 10854 25834 10906
rect 25846 10854 25898 10906
rect 25910 10854 25962 10906
rect 25974 10854 26026 10906
rect 8116 10752 8168 10804
rect 11152 10752 11204 10804
rect 11612 10752 11664 10804
rect 13544 10752 13596 10804
rect 17684 10795 17736 10804
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 17776 10752 17828 10804
rect 19432 10795 19484 10804
rect 19432 10761 19441 10795
rect 19441 10761 19475 10795
rect 19475 10761 19484 10795
rect 19432 10752 19484 10761
rect 19616 10752 19668 10804
rect 12624 10727 12676 10736
rect 12624 10693 12633 10727
rect 12633 10693 12667 10727
rect 12667 10693 12676 10727
rect 12624 10684 12676 10693
rect 14556 10684 14608 10736
rect 15476 10684 15528 10736
rect 17316 10727 17368 10736
rect 17316 10693 17325 10727
rect 17325 10693 17359 10727
rect 17359 10693 17368 10727
rect 17316 10684 17368 10693
rect 19248 10684 19300 10736
rect 22284 10752 22336 10804
rect 6736 10412 6788 10464
rect 8944 10659 8996 10668
rect 8300 10591 8352 10600
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 8300 10548 8352 10557
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9036 10616 9088 10668
rect 10324 10616 10376 10668
rect 11888 10616 11940 10668
rect 13544 10616 13596 10668
rect 18880 10659 18932 10668
rect 14740 10548 14792 10600
rect 16212 10548 16264 10600
rect 16304 10548 16356 10600
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 20904 10659 20956 10668
rect 20904 10625 20913 10659
rect 20913 10625 20947 10659
rect 20947 10625 20956 10659
rect 20904 10616 20956 10625
rect 21732 10616 21784 10668
rect 18972 10548 19024 10600
rect 20076 10548 20128 10600
rect 20996 10548 21048 10600
rect 21916 10548 21968 10600
rect 7656 10412 7708 10464
rect 9128 10480 9180 10532
rect 11152 10480 11204 10532
rect 23848 10480 23900 10532
rect 8300 10412 8352 10464
rect 9588 10412 9640 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12992 10412 13044 10464
rect 13820 10412 13872 10464
rect 15844 10412 15896 10464
rect 21640 10412 21692 10464
rect 22192 10455 22244 10464
rect 22192 10421 22201 10455
rect 22201 10421 22235 10455
rect 22235 10421 22244 10455
rect 22192 10412 22244 10421
rect 22468 10455 22520 10464
rect 22468 10421 22477 10455
rect 22477 10421 22511 10455
rect 22511 10421 22520 10455
rect 22468 10412 22520 10421
rect 3282 10310 3334 10362
rect 3346 10310 3398 10362
rect 3410 10310 3462 10362
rect 3474 10310 3526 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 6410 10310 6462 10362
rect 6474 10310 6526 10362
rect 9282 10310 9334 10362
rect 9346 10310 9398 10362
rect 9410 10310 9462 10362
rect 9474 10310 9526 10362
rect 12282 10310 12334 10362
rect 12346 10310 12398 10362
rect 12410 10310 12462 10362
rect 12474 10310 12526 10362
rect 15282 10310 15334 10362
rect 15346 10310 15398 10362
rect 15410 10310 15462 10362
rect 15474 10310 15526 10362
rect 18282 10310 18334 10362
rect 18346 10310 18398 10362
rect 18410 10310 18462 10362
rect 18474 10310 18526 10362
rect 21282 10310 21334 10362
rect 21346 10310 21398 10362
rect 21410 10310 21462 10362
rect 21474 10310 21526 10362
rect 24282 10310 24334 10362
rect 24346 10310 24398 10362
rect 24410 10310 24462 10362
rect 24474 10310 24526 10362
rect 27282 10310 27334 10362
rect 27346 10310 27398 10362
rect 27410 10310 27462 10362
rect 27474 10310 27526 10362
rect 6736 10208 6788 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 10692 10208 10744 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 14556 10208 14608 10260
rect 14740 10208 14792 10260
rect 14832 10208 14884 10260
rect 8300 10140 8352 10192
rect 11980 10140 12032 10192
rect 10416 10115 10468 10124
rect 6184 10047 6236 10056
rect 6184 10013 6193 10047
rect 6193 10013 6227 10047
rect 6227 10013 6236 10047
rect 6184 10004 6236 10013
rect 6920 10004 6972 10056
rect 10416 10081 10425 10115
rect 10425 10081 10459 10115
rect 10459 10081 10468 10115
rect 10416 10072 10468 10081
rect 13820 10072 13872 10124
rect 16212 10072 16264 10124
rect 8300 10047 8352 10056
rect 7288 9936 7340 9988
rect 7564 9936 7616 9988
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 13360 10004 13412 10056
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 16672 10208 16724 10260
rect 19524 10208 19576 10260
rect 21180 10208 21232 10260
rect 20536 10140 20588 10192
rect 20904 10140 20956 10192
rect 20076 10072 20128 10124
rect 20720 10072 20772 10124
rect 22100 10072 22152 10124
rect 23848 10115 23900 10124
rect 23848 10081 23857 10115
rect 23857 10081 23891 10115
rect 23891 10081 23900 10115
rect 23848 10072 23900 10081
rect 19524 10004 19576 10056
rect 10600 9936 10652 9988
rect 11152 9936 11204 9988
rect 12164 9936 12216 9988
rect 16028 9979 16080 9988
rect 10324 9868 10376 9920
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 15384 9868 15436 9920
rect 16028 9945 16037 9979
rect 16037 9945 16071 9979
rect 16071 9945 16080 9979
rect 16028 9936 16080 9945
rect 16672 9979 16724 9988
rect 16672 9945 16681 9979
rect 16681 9945 16715 9979
rect 16715 9945 16724 9979
rect 16672 9936 16724 9945
rect 18696 9979 18748 9988
rect 18696 9945 18705 9979
rect 18705 9945 18739 9979
rect 18739 9945 18748 9979
rect 18696 9936 18748 9945
rect 22100 9979 22152 9988
rect 22100 9945 22109 9979
rect 22109 9945 22143 9979
rect 22143 9945 22152 9979
rect 22100 9936 22152 9945
rect 19064 9868 19116 9920
rect 20076 9868 20128 9920
rect 22008 9868 22060 9920
rect 1782 9766 1834 9818
rect 1846 9766 1898 9818
rect 1910 9766 1962 9818
rect 1974 9766 2026 9818
rect 4782 9766 4834 9818
rect 4846 9766 4898 9818
rect 4910 9766 4962 9818
rect 4974 9766 5026 9818
rect 7782 9766 7834 9818
rect 7846 9766 7898 9818
rect 7910 9766 7962 9818
rect 7974 9766 8026 9818
rect 10782 9766 10834 9818
rect 10846 9766 10898 9818
rect 10910 9766 10962 9818
rect 10974 9766 11026 9818
rect 13782 9766 13834 9818
rect 13846 9766 13898 9818
rect 13910 9766 13962 9818
rect 13974 9766 14026 9818
rect 16782 9766 16834 9818
rect 16846 9766 16898 9818
rect 16910 9766 16962 9818
rect 16974 9766 17026 9818
rect 19782 9766 19834 9818
rect 19846 9766 19898 9818
rect 19910 9766 19962 9818
rect 19974 9766 20026 9818
rect 22782 9766 22834 9818
rect 22846 9766 22898 9818
rect 22910 9766 22962 9818
rect 22974 9766 23026 9818
rect 25782 9766 25834 9818
rect 25846 9766 25898 9818
rect 25910 9766 25962 9818
rect 25974 9766 26026 9818
rect 8300 9664 8352 9716
rect 8668 9664 8720 9716
rect 10416 9664 10468 9716
rect 11152 9664 11204 9716
rect 11888 9664 11940 9716
rect 13636 9664 13688 9716
rect 6184 9596 6236 9648
rect 7564 9596 7616 9648
rect 7748 9596 7800 9648
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 11244 9596 11296 9648
rect 13360 9596 13412 9648
rect 14924 9664 14976 9716
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 22008 9707 22060 9716
rect 22008 9673 22017 9707
rect 22017 9673 22051 9707
rect 22051 9673 22060 9707
rect 22008 9664 22060 9673
rect 22100 9664 22152 9716
rect 16304 9596 16356 9648
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 9588 9460 9640 9512
rect 10600 9460 10652 9512
rect 11520 9528 11572 9580
rect 11888 9528 11940 9580
rect 14464 9528 14516 9580
rect 16120 9528 16172 9580
rect 16580 9528 16632 9580
rect 17500 9596 17552 9648
rect 21088 9596 21140 9648
rect 19064 9571 19116 9580
rect 10784 9460 10836 9512
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 9128 9392 9180 9444
rect 13544 9460 13596 9512
rect 14188 9460 14240 9512
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 19064 9537 19073 9571
rect 19073 9537 19107 9571
rect 19107 9537 19116 9571
rect 19064 9528 19116 9537
rect 19248 9571 19300 9580
rect 19248 9537 19257 9571
rect 19257 9537 19291 9571
rect 19291 9537 19300 9571
rect 19248 9528 19300 9537
rect 19524 9528 19576 9580
rect 21824 9571 21876 9580
rect 21824 9537 21833 9571
rect 21833 9537 21867 9571
rect 21867 9537 21876 9571
rect 21824 9528 21876 9537
rect 21916 9528 21968 9580
rect 18972 9460 19024 9512
rect 19984 9392 20036 9444
rect 22284 9503 22336 9512
rect 22284 9469 22293 9503
rect 22293 9469 22327 9503
rect 22327 9469 22336 9503
rect 22284 9460 22336 9469
rect 20536 9435 20588 9444
rect 20536 9401 20545 9435
rect 20545 9401 20579 9435
rect 20579 9401 20588 9435
rect 20536 9392 20588 9401
rect 21088 9392 21140 9444
rect 22192 9392 22244 9444
rect 13360 9324 13412 9376
rect 14188 9324 14240 9376
rect 17132 9324 17184 9376
rect 20076 9324 20128 9376
rect 21732 9324 21784 9376
rect 3282 9222 3334 9274
rect 3346 9222 3398 9274
rect 3410 9222 3462 9274
rect 3474 9222 3526 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 6410 9222 6462 9274
rect 6474 9222 6526 9274
rect 9282 9222 9334 9274
rect 9346 9222 9398 9274
rect 9410 9222 9462 9274
rect 9474 9222 9526 9274
rect 12282 9222 12334 9274
rect 12346 9222 12398 9274
rect 12410 9222 12462 9274
rect 12474 9222 12526 9274
rect 15282 9222 15334 9274
rect 15346 9222 15398 9274
rect 15410 9222 15462 9274
rect 15474 9222 15526 9274
rect 18282 9222 18334 9274
rect 18346 9222 18398 9274
rect 18410 9222 18462 9274
rect 18474 9222 18526 9274
rect 21282 9222 21334 9274
rect 21346 9222 21398 9274
rect 21410 9222 21462 9274
rect 21474 9222 21526 9274
rect 24282 9222 24334 9274
rect 24346 9222 24398 9274
rect 24410 9222 24462 9274
rect 24474 9222 24526 9274
rect 27282 9222 27334 9274
rect 27346 9222 27398 9274
rect 27410 9222 27462 9274
rect 27474 9222 27526 9274
rect 7288 9120 7340 9172
rect 8300 9120 8352 9172
rect 9128 9120 9180 9172
rect 10600 9120 10652 9172
rect 10784 9120 10836 9172
rect 16120 9163 16172 9172
rect 16120 9129 16129 9163
rect 16129 9129 16163 9163
rect 16163 9129 16172 9163
rect 16120 9120 16172 9129
rect 16580 9163 16632 9172
rect 16580 9129 16589 9163
rect 16589 9129 16623 9163
rect 16623 9129 16632 9163
rect 16580 9120 16632 9129
rect 18696 9120 18748 9172
rect 19248 9120 19300 9172
rect 22100 9120 22152 9172
rect 7748 9052 7800 9104
rect 21916 9052 21968 9104
rect 6736 8984 6788 9036
rect 7104 8984 7156 9036
rect 8668 8984 8720 9036
rect 10508 8984 10560 9036
rect 13452 8984 13504 9036
rect 15844 8984 15896 9036
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 18880 9027 18932 9036
rect 18880 8993 18889 9027
rect 18889 8993 18923 9027
rect 18923 8993 18932 9027
rect 18880 8984 18932 8993
rect 21088 9027 21140 9036
rect 21088 8993 21097 9027
rect 21097 8993 21131 9027
rect 21131 8993 21140 9027
rect 21088 8984 21140 8993
rect 6092 8916 6144 8968
rect 8116 8916 8168 8968
rect 9864 8891 9916 8900
rect 9864 8857 9873 8891
rect 9873 8857 9907 8891
rect 9907 8857 9916 8891
rect 9864 8848 9916 8857
rect 10140 8916 10192 8968
rect 12164 8916 12216 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 10232 8848 10284 8900
rect 11796 8848 11848 8900
rect 13176 8848 13228 8900
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 16672 8916 16724 8968
rect 19156 8916 19208 8968
rect 19984 8916 20036 8968
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 21640 8916 21692 8968
rect 22284 8916 22336 8968
rect 17684 8848 17736 8900
rect 19340 8848 19392 8900
rect 20720 8848 20772 8900
rect 22192 8848 22244 8900
rect 14464 8780 14516 8832
rect 20076 8780 20128 8832
rect 1782 8678 1834 8730
rect 1846 8678 1898 8730
rect 1910 8678 1962 8730
rect 1974 8678 2026 8730
rect 4782 8678 4834 8730
rect 4846 8678 4898 8730
rect 4910 8678 4962 8730
rect 4974 8678 5026 8730
rect 7782 8678 7834 8730
rect 7846 8678 7898 8730
rect 7910 8678 7962 8730
rect 7974 8678 8026 8730
rect 10782 8678 10834 8730
rect 10846 8678 10898 8730
rect 10910 8678 10962 8730
rect 10974 8678 11026 8730
rect 13782 8678 13834 8730
rect 13846 8678 13898 8730
rect 13910 8678 13962 8730
rect 13974 8678 14026 8730
rect 16782 8678 16834 8730
rect 16846 8678 16898 8730
rect 16910 8678 16962 8730
rect 16974 8678 17026 8730
rect 19782 8678 19834 8730
rect 19846 8678 19898 8730
rect 19910 8678 19962 8730
rect 19974 8678 20026 8730
rect 22782 8678 22834 8730
rect 22846 8678 22898 8730
rect 22910 8678 22962 8730
rect 22974 8678 23026 8730
rect 25782 8678 25834 8730
rect 25846 8678 25898 8730
rect 25910 8678 25962 8730
rect 25974 8678 26026 8730
rect 7380 8576 7432 8628
rect 8116 8576 8168 8628
rect 8760 8576 8812 8628
rect 11520 8576 11572 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 13360 8576 13412 8628
rect 16672 8576 16724 8628
rect 17132 8576 17184 8628
rect 17684 8619 17736 8628
rect 17684 8585 17693 8619
rect 17693 8585 17727 8619
rect 17727 8585 17736 8619
rect 17684 8576 17736 8585
rect 18604 8576 18656 8628
rect 18788 8576 18840 8628
rect 19156 8576 19208 8628
rect 20536 8576 20588 8628
rect 21180 8619 21232 8628
rect 21180 8585 21189 8619
rect 21189 8585 21223 8619
rect 21223 8585 21232 8619
rect 21180 8576 21232 8585
rect 21272 8576 21324 8628
rect 21824 8576 21876 8628
rect 22192 8576 22244 8628
rect 7656 8551 7708 8560
rect 7656 8517 7665 8551
rect 7665 8517 7699 8551
rect 7699 8517 7708 8551
rect 7656 8508 7708 8517
rect 8576 8508 8628 8560
rect 8300 8440 8352 8492
rect 10048 8508 10100 8560
rect 13636 8508 13688 8560
rect 14464 8508 14516 8560
rect 15660 8508 15712 8560
rect 11428 8483 11480 8492
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 9588 8372 9640 8424
rect 10784 8415 10836 8424
rect 10784 8381 10793 8415
rect 10793 8381 10827 8415
rect 10827 8381 10836 8415
rect 10784 8372 10836 8381
rect 11428 8449 11437 8483
rect 11437 8449 11471 8483
rect 11471 8449 11480 8483
rect 11428 8440 11480 8449
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 17776 8440 17828 8492
rect 18880 8440 18932 8492
rect 11244 8372 11296 8424
rect 11980 8372 12032 8424
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 7564 8304 7616 8356
rect 11152 8304 11204 8356
rect 16672 8304 16724 8356
rect 19340 8304 19392 8356
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19708 8483 19760 8492
rect 19524 8440 19576 8449
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 19708 8440 19760 8449
rect 20444 8508 20496 8560
rect 22008 8508 22060 8560
rect 20076 8304 20128 8356
rect 21640 8440 21692 8492
rect 20628 8415 20680 8424
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 6092 8236 6144 8288
rect 14556 8236 14608 8288
rect 16304 8236 16356 8288
rect 19248 8236 19300 8288
rect 22468 8304 22520 8356
rect 22284 8279 22336 8288
rect 22284 8245 22293 8279
rect 22293 8245 22327 8279
rect 22327 8245 22336 8279
rect 22284 8236 22336 8245
rect 3282 8134 3334 8186
rect 3346 8134 3398 8186
rect 3410 8134 3462 8186
rect 3474 8134 3526 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 6410 8134 6462 8186
rect 6474 8134 6526 8186
rect 9282 8134 9334 8186
rect 9346 8134 9398 8186
rect 9410 8134 9462 8186
rect 9474 8134 9526 8186
rect 12282 8134 12334 8186
rect 12346 8134 12398 8186
rect 12410 8134 12462 8186
rect 12474 8134 12526 8186
rect 15282 8134 15334 8186
rect 15346 8134 15398 8186
rect 15410 8134 15462 8186
rect 15474 8134 15526 8186
rect 18282 8134 18334 8186
rect 18346 8134 18398 8186
rect 18410 8134 18462 8186
rect 18474 8134 18526 8186
rect 21282 8134 21334 8186
rect 21346 8134 21398 8186
rect 21410 8134 21462 8186
rect 21474 8134 21526 8186
rect 24282 8134 24334 8186
rect 24346 8134 24398 8186
rect 24410 8134 24462 8186
rect 24474 8134 24526 8186
rect 27282 8134 27334 8186
rect 27346 8134 27398 8186
rect 27410 8134 27462 8186
rect 27474 8134 27526 8186
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 9036 8075 9088 8084
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 9128 8032 9180 8084
rect 10232 8032 10284 8084
rect 13176 8032 13228 8084
rect 13452 8032 13504 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 16212 8075 16264 8084
rect 16212 8041 16221 8075
rect 16221 8041 16255 8075
rect 16255 8041 16264 8075
rect 16212 8032 16264 8041
rect 19064 8032 19116 8084
rect 22284 8032 22336 8084
rect 8760 7964 8812 8016
rect 10140 7964 10192 8016
rect 11428 7964 11480 8016
rect 19708 8007 19760 8016
rect 19708 7973 19717 8007
rect 19717 7973 19751 8007
rect 19751 7973 19760 8007
rect 19708 7964 19760 7973
rect 20812 7964 20864 8016
rect 8300 7939 8352 7948
rect 8300 7905 8309 7939
rect 8309 7905 8343 7939
rect 8343 7905 8352 7939
rect 8300 7896 8352 7905
rect 10784 7896 10836 7948
rect 13544 7896 13596 7948
rect 16028 7896 16080 7948
rect 6184 7828 6236 7880
rect 7012 7828 7064 7880
rect 8760 7871 8812 7880
rect 7472 7760 7524 7812
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 9588 7828 9640 7880
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 10140 7871 10192 7880
rect 9956 7828 10008 7837
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10324 7828 10376 7880
rect 13360 7871 13412 7880
rect 10232 7760 10284 7812
rect 12716 7760 12768 7812
rect 11520 7692 11572 7744
rect 12256 7735 12308 7744
rect 12256 7701 12265 7735
rect 12265 7701 12299 7735
rect 12299 7701 12308 7735
rect 12256 7692 12308 7701
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 19156 7896 19208 7948
rect 22008 7939 22060 7948
rect 22008 7905 22017 7939
rect 22017 7905 22051 7939
rect 22051 7905 22060 7939
rect 22008 7896 22060 7905
rect 18236 7828 18288 7880
rect 19524 7828 19576 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 18696 7760 18748 7812
rect 21180 7760 21232 7812
rect 13636 7692 13688 7744
rect 16304 7692 16356 7744
rect 19248 7692 19300 7744
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 1782 7590 1834 7642
rect 1846 7590 1898 7642
rect 1910 7590 1962 7642
rect 1974 7590 2026 7642
rect 4782 7590 4834 7642
rect 4846 7590 4898 7642
rect 4910 7590 4962 7642
rect 4974 7590 5026 7642
rect 7782 7590 7834 7642
rect 7846 7590 7898 7642
rect 7910 7590 7962 7642
rect 7974 7590 8026 7642
rect 10782 7590 10834 7642
rect 10846 7590 10898 7642
rect 10910 7590 10962 7642
rect 10974 7590 11026 7642
rect 13782 7590 13834 7642
rect 13846 7590 13898 7642
rect 13910 7590 13962 7642
rect 13974 7590 14026 7642
rect 16782 7590 16834 7642
rect 16846 7590 16898 7642
rect 16910 7590 16962 7642
rect 16974 7590 17026 7642
rect 19782 7590 19834 7642
rect 19846 7590 19898 7642
rect 19910 7590 19962 7642
rect 19974 7590 20026 7642
rect 22782 7590 22834 7642
rect 22846 7590 22898 7642
rect 22910 7590 22962 7642
rect 22974 7590 23026 7642
rect 25782 7590 25834 7642
rect 25846 7590 25898 7642
rect 25910 7590 25962 7642
rect 25974 7590 26026 7642
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 8300 7488 8352 7540
rect 9864 7488 9916 7540
rect 10232 7488 10284 7540
rect 13360 7488 13412 7540
rect 16672 7531 16724 7540
rect 16672 7497 16681 7531
rect 16681 7497 16715 7531
rect 16715 7497 16724 7531
rect 16672 7488 16724 7497
rect 17776 7488 17828 7540
rect 18236 7531 18288 7540
rect 18236 7497 18245 7531
rect 18245 7497 18279 7531
rect 18279 7497 18288 7531
rect 18236 7488 18288 7497
rect 20444 7531 20496 7540
rect 20444 7497 20453 7531
rect 20453 7497 20487 7531
rect 20487 7497 20496 7531
rect 20444 7488 20496 7497
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 21732 7488 21784 7540
rect 7104 7420 7156 7472
rect 9956 7420 10008 7472
rect 10140 7420 10192 7472
rect 11520 7420 11572 7472
rect 12256 7420 12308 7472
rect 12900 7420 12952 7472
rect 14556 7420 14608 7472
rect 21180 7463 21232 7472
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 13268 7395 13320 7404
rect 6092 7284 6144 7336
rect 10324 7284 10376 7336
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 13544 7352 13596 7404
rect 14740 7395 14792 7404
rect 10876 7284 10928 7336
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 21180 7429 21189 7463
rect 21189 7429 21223 7463
rect 21223 7429 21232 7463
rect 21180 7420 21232 7429
rect 14832 7352 14884 7361
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 16120 7352 16172 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 22008 7352 22060 7404
rect 19340 7327 19392 7336
rect 19340 7293 19349 7327
rect 19349 7293 19383 7327
rect 19383 7293 19392 7327
rect 19340 7284 19392 7293
rect 21732 7284 21784 7336
rect 10048 7148 10100 7200
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 11152 7148 11204 7200
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12072 7148 12124 7157
rect 14280 7216 14332 7268
rect 14924 7216 14976 7268
rect 19248 7216 19300 7268
rect 14372 7148 14424 7200
rect 16120 7148 16172 7200
rect 18972 7148 19024 7200
rect 19616 7148 19668 7200
rect 3282 7046 3334 7098
rect 3346 7046 3398 7098
rect 3410 7046 3462 7098
rect 3474 7046 3526 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 6410 7046 6462 7098
rect 6474 7046 6526 7098
rect 9282 7046 9334 7098
rect 9346 7046 9398 7098
rect 9410 7046 9462 7098
rect 9474 7046 9526 7098
rect 12282 7046 12334 7098
rect 12346 7046 12398 7098
rect 12410 7046 12462 7098
rect 12474 7046 12526 7098
rect 15282 7046 15334 7098
rect 15346 7046 15398 7098
rect 15410 7046 15462 7098
rect 15474 7046 15526 7098
rect 18282 7046 18334 7098
rect 18346 7046 18398 7098
rect 18410 7046 18462 7098
rect 18474 7046 18526 7098
rect 21282 7046 21334 7098
rect 21346 7046 21398 7098
rect 21410 7046 21462 7098
rect 21474 7046 21526 7098
rect 24282 7046 24334 7098
rect 24346 7046 24398 7098
rect 24410 7046 24462 7098
rect 24474 7046 24526 7098
rect 27282 7046 27334 7098
rect 27346 7046 27398 7098
rect 27410 7046 27462 7098
rect 27474 7046 27526 7098
rect 9864 6944 9916 6996
rect 10876 6987 10928 6996
rect 10876 6953 10885 6987
rect 10885 6953 10919 6987
rect 10919 6953 10928 6987
rect 10876 6944 10928 6953
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 9128 6876 9180 6928
rect 11796 6944 11848 6996
rect 13268 6944 13320 6996
rect 14556 6987 14608 6996
rect 14556 6953 14565 6987
rect 14565 6953 14599 6987
rect 14599 6953 14608 6987
rect 14556 6944 14608 6953
rect 14740 6944 14792 6996
rect 16304 6987 16356 6996
rect 16304 6953 16313 6987
rect 16313 6953 16347 6987
rect 16347 6953 16356 6987
rect 16304 6944 16356 6953
rect 16672 6944 16724 6996
rect 17684 6944 17736 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 15108 6876 15160 6928
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 14832 6808 14884 6860
rect 15660 6808 15712 6860
rect 20076 6808 20128 6860
rect 10048 6783 10100 6792
rect 6828 6672 6880 6724
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 15844 6740 15896 6792
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 19432 6740 19484 6792
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 12164 6672 12216 6724
rect 15936 6672 15988 6724
rect 6644 6604 6696 6656
rect 17960 6604 18012 6656
rect 19340 6604 19392 6656
rect 21180 6740 21232 6792
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 20168 6604 20220 6656
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 22008 6604 22060 6656
rect 1782 6502 1834 6554
rect 1846 6502 1898 6554
rect 1910 6502 1962 6554
rect 1974 6502 2026 6554
rect 4782 6502 4834 6554
rect 4846 6502 4898 6554
rect 4910 6502 4962 6554
rect 4974 6502 5026 6554
rect 7782 6502 7834 6554
rect 7846 6502 7898 6554
rect 7910 6502 7962 6554
rect 7974 6502 8026 6554
rect 10782 6502 10834 6554
rect 10846 6502 10898 6554
rect 10910 6502 10962 6554
rect 10974 6502 11026 6554
rect 13782 6502 13834 6554
rect 13846 6502 13898 6554
rect 13910 6502 13962 6554
rect 13974 6502 14026 6554
rect 16782 6502 16834 6554
rect 16846 6502 16898 6554
rect 16910 6502 16962 6554
rect 16974 6502 17026 6554
rect 19782 6502 19834 6554
rect 19846 6502 19898 6554
rect 19910 6502 19962 6554
rect 19974 6502 20026 6554
rect 22782 6502 22834 6554
rect 22846 6502 22898 6554
rect 22910 6502 22962 6554
rect 22974 6502 23026 6554
rect 25782 6502 25834 6554
rect 25846 6502 25898 6554
rect 25910 6502 25962 6554
rect 25974 6502 26026 6554
rect 7472 6400 7524 6452
rect 9588 6400 9640 6452
rect 10048 6400 10100 6452
rect 10600 6400 10652 6452
rect 12164 6400 12216 6452
rect 12716 6400 12768 6452
rect 15844 6400 15896 6452
rect 5356 6375 5408 6384
rect 5356 6341 5365 6375
rect 5365 6341 5399 6375
rect 5399 6341 5408 6375
rect 5356 6332 5408 6341
rect 9864 6332 9916 6384
rect 11704 6332 11756 6384
rect 15660 6375 15712 6384
rect 15660 6341 15669 6375
rect 15669 6341 15703 6375
rect 15703 6341 15712 6375
rect 15660 6332 15712 6341
rect 18880 6332 18932 6384
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 6276 6307 6328 6316
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 7656 6264 7708 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 9956 6307 10008 6316
rect 8760 6264 8812 6273
rect 7012 6196 7064 6248
rect 8668 6196 8720 6248
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 11336 6307 11388 6316
rect 11336 6273 11345 6307
rect 11345 6273 11379 6307
rect 11379 6273 11388 6307
rect 11336 6264 11388 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 14648 6264 14700 6316
rect 15936 6264 15988 6316
rect 21640 6332 21692 6384
rect 19524 6264 19576 6316
rect 20628 6264 20680 6316
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 16580 6196 16632 6248
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 19616 6239 19668 6248
rect 8300 6128 8352 6180
rect 18788 6128 18840 6180
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 20996 6239 21048 6248
rect 20996 6205 21005 6239
rect 21005 6205 21039 6239
rect 21039 6205 21048 6239
rect 20996 6196 21048 6205
rect 22008 6196 22060 6248
rect 20076 6128 20128 6180
rect 14464 6060 14516 6112
rect 16672 6060 16724 6112
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 3282 5958 3334 6010
rect 3346 5958 3398 6010
rect 3410 5958 3462 6010
rect 3474 5958 3526 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 6410 5958 6462 6010
rect 6474 5958 6526 6010
rect 9282 5958 9334 6010
rect 9346 5958 9398 6010
rect 9410 5958 9462 6010
rect 9474 5958 9526 6010
rect 12282 5958 12334 6010
rect 12346 5958 12398 6010
rect 12410 5958 12462 6010
rect 12474 5958 12526 6010
rect 15282 5958 15334 6010
rect 15346 5958 15398 6010
rect 15410 5958 15462 6010
rect 15474 5958 15526 6010
rect 18282 5958 18334 6010
rect 18346 5958 18398 6010
rect 18410 5958 18462 6010
rect 18474 5958 18526 6010
rect 21282 5958 21334 6010
rect 21346 5958 21398 6010
rect 21410 5958 21462 6010
rect 21474 5958 21526 6010
rect 24282 5958 24334 6010
rect 24346 5958 24398 6010
rect 24410 5958 24462 6010
rect 24474 5958 24526 6010
rect 27282 5958 27334 6010
rect 27346 5958 27398 6010
rect 27410 5958 27462 6010
rect 27474 5958 27526 6010
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 5540 5856 5592 5908
rect 6828 5856 6880 5908
rect 7656 5856 7708 5908
rect 11336 5856 11388 5908
rect 12992 5788 13044 5840
rect 17960 5831 18012 5840
rect 6736 5763 6788 5772
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 7012 5763 7064 5772
rect 7012 5729 7021 5763
rect 7021 5729 7055 5763
rect 7055 5729 7064 5763
rect 7012 5720 7064 5729
rect 9128 5720 9180 5772
rect 13084 5720 13136 5772
rect 14464 5720 14516 5772
rect 16212 5720 16264 5772
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 12808 5695 12860 5704
rect 9956 5652 10008 5661
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 12992 5652 13044 5704
rect 14280 5652 14332 5704
rect 15936 5652 15988 5704
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 17960 5797 17969 5831
rect 17969 5797 18003 5831
rect 18003 5797 18012 5831
rect 17960 5788 18012 5797
rect 19524 5856 19576 5908
rect 20720 5856 20772 5908
rect 21180 5788 21232 5840
rect 18788 5763 18840 5772
rect 18788 5729 18797 5763
rect 18797 5729 18831 5763
rect 18831 5729 18840 5763
rect 18788 5720 18840 5729
rect 20996 5720 21048 5772
rect 21824 5763 21876 5772
rect 21824 5729 21833 5763
rect 21833 5729 21867 5763
rect 21867 5729 21876 5763
rect 21824 5720 21876 5729
rect 22008 5763 22060 5772
rect 22008 5729 22017 5763
rect 22017 5729 22051 5763
rect 22051 5729 22060 5763
rect 22008 5720 22060 5729
rect 16488 5652 16540 5661
rect 17132 5652 17184 5704
rect 17960 5652 18012 5704
rect 18604 5652 18656 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 21732 5695 21784 5704
rect 21732 5661 21741 5695
rect 21741 5661 21775 5695
rect 21775 5661 21784 5695
rect 21732 5652 21784 5661
rect 6644 5584 6696 5636
rect 11244 5627 11296 5636
rect 11244 5593 11253 5627
rect 11253 5593 11287 5627
rect 11287 5593 11296 5627
rect 11244 5584 11296 5593
rect 11428 5627 11480 5636
rect 11428 5593 11437 5627
rect 11437 5593 11471 5627
rect 11471 5593 11480 5627
rect 11428 5584 11480 5593
rect 11612 5627 11664 5636
rect 11612 5593 11621 5627
rect 11621 5593 11655 5627
rect 11655 5593 11664 5627
rect 11612 5584 11664 5593
rect 8668 5516 8720 5568
rect 11520 5559 11572 5568
rect 11520 5525 11529 5559
rect 11529 5525 11563 5559
rect 11563 5525 11572 5559
rect 16028 5584 16080 5636
rect 21364 5584 21416 5636
rect 11520 5516 11572 5525
rect 13544 5516 13596 5568
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 16580 5516 16632 5568
rect 1782 5414 1834 5466
rect 1846 5414 1898 5466
rect 1910 5414 1962 5466
rect 1974 5414 2026 5466
rect 4782 5414 4834 5466
rect 4846 5414 4898 5466
rect 4910 5414 4962 5466
rect 4974 5414 5026 5466
rect 7782 5414 7834 5466
rect 7846 5414 7898 5466
rect 7910 5414 7962 5466
rect 7974 5414 8026 5466
rect 10782 5414 10834 5466
rect 10846 5414 10898 5466
rect 10910 5414 10962 5466
rect 10974 5414 11026 5466
rect 13782 5414 13834 5466
rect 13846 5414 13898 5466
rect 13910 5414 13962 5466
rect 13974 5414 14026 5466
rect 16782 5414 16834 5466
rect 16846 5414 16898 5466
rect 16910 5414 16962 5466
rect 16974 5414 17026 5466
rect 19782 5414 19834 5466
rect 19846 5414 19898 5466
rect 19910 5414 19962 5466
rect 19974 5414 20026 5466
rect 22782 5414 22834 5466
rect 22846 5414 22898 5466
rect 22910 5414 22962 5466
rect 22974 5414 23026 5466
rect 25782 5414 25834 5466
rect 25846 5414 25898 5466
rect 25910 5414 25962 5466
rect 25974 5414 26026 5466
rect 6644 5312 6696 5364
rect 7012 5312 7064 5364
rect 8116 5355 8168 5364
rect 8116 5321 8125 5355
rect 8125 5321 8159 5355
rect 8159 5321 8168 5355
rect 8116 5312 8168 5321
rect 15936 5312 15988 5364
rect 18604 5312 18656 5364
rect 21640 5312 21692 5364
rect 21824 5355 21876 5364
rect 21824 5321 21833 5355
rect 21833 5321 21867 5355
rect 21867 5321 21876 5355
rect 21824 5312 21876 5321
rect 8300 5244 8352 5296
rect 8668 5287 8720 5296
rect 8668 5253 8677 5287
rect 8677 5253 8711 5287
rect 8711 5253 8720 5287
rect 8668 5244 8720 5253
rect 9128 5244 9180 5296
rect 11612 5287 11664 5296
rect 6736 5176 6788 5228
rect 9588 5176 9640 5228
rect 11612 5253 11621 5287
rect 11621 5253 11655 5287
rect 11655 5253 11664 5287
rect 11612 5244 11664 5253
rect 14924 5244 14976 5296
rect 16672 5287 16724 5296
rect 16672 5253 16681 5287
rect 16681 5253 16715 5287
rect 16715 5253 16724 5287
rect 16672 5244 16724 5253
rect 18972 5287 19024 5296
rect 18972 5253 18981 5287
rect 18981 5253 19015 5287
rect 19015 5253 19024 5287
rect 18972 5244 19024 5253
rect 19708 5244 19760 5296
rect 21364 5287 21416 5296
rect 21364 5253 21373 5287
rect 21373 5253 21407 5287
rect 21407 5253 21416 5287
rect 21364 5244 21416 5253
rect 11152 5219 11204 5228
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 11428 5176 11480 5228
rect 11888 5176 11940 5228
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 14648 5219 14700 5228
rect 14648 5185 14657 5219
rect 14657 5185 14691 5219
rect 14691 5185 14700 5219
rect 14648 5176 14700 5185
rect 16212 5219 16264 5228
rect 16212 5185 16241 5219
rect 16241 5185 16264 5219
rect 16212 5176 16264 5185
rect 12716 5151 12768 5160
rect 9128 5040 9180 5092
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 12992 5108 13044 5160
rect 14372 5108 14424 5160
rect 17776 5108 17828 5160
rect 19064 5108 19116 5160
rect 20168 5108 20220 5160
rect 11244 5040 11296 5092
rect 18604 5040 18656 5092
rect 10232 5015 10284 5024
rect 10232 4981 10241 5015
rect 10241 4981 10275 5015
rect 10275 4981 10284 5015
rect 10232 4972 10284 4981
rect 14740 4972 14792 5024
rect 16488 4972 16540 5024
rect 3282 4870 3334 4922
rect 3346 4870 3398 4922
rect 3410 4870 3462 4922
rect 3474 4870 3526 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 6410 4870 6462 4922
rect 6474 4870 6526 4922
rect 9282 4870 9334 4922
rect 9346 4870 9398 4922
rect 9410 4870 9462 4922
rect 9474 4870 9526 4922
rect 12282 4870 12334 4922
rect 12346 4870 12398 4922
rect 12410 4870 12462 4922
rect 12474 4870 12526 4922
rect 15282 4870 15334 4922
rect 15346 4870 15398 4922
rect 15410 4870 15462 4922
rect 15474 4870 15526 4922
rect 18282 4870 18334 4922
rect 18346 4870 18398 4922
rect 18410 4870 18462 4922
rect 18474 4870 18526 4922
rect 21282 4870 21334 4922
rect 21346 4870 21398 4922
rect 21410 4870 21462 4922
rect 21474 4870 21526 4922
rect 24282 4870 24334 4922
rect 24346 4870 24398 4922
rect 24410 4870 24462 4922
rect 24474 4870 24526 4922
rect 27282 4870 27334 4922
rect 27346 4870 27398 4922
rect 27410 4870 27462 4922
rect 27474 4870 27526 4922
rect 6828 4811 6880 4820
rect 6828 4777 6837 4811
rect 6837 4777 6871 4811
rect 6871 4777 6880 4811
rect 6828 4768 6880 4777
rect 8760 4768 8812 4820
rect 9128 4811 9180 4820
rect 9128 4777 9137 4811
rect 9137 4777 9171 4811
rect 9171 4777 9180 4811
rect 9128 4768 9180 4777
rect 11888 4811 11940 4820
rect 11888 4777 11897 4811
rect 11897 4777 11931 4811
rect 11931 4777 11940 4811
rect 11888 4768 11940 4777
rect 14464 4768 14516 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 18972 4768 19024 4820
rect 19708 4768 19760 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 22008 4768 22060 4820
rect 18604 4700 18656 4752
rect 19064 4700 19116 4752
rect 20720 4700 20772 4752
rect 21732 4700 21784 4752
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 6644 4428 6696 4480
rect 8300 4564 8352 4616
rect 9588 4564 9640 4616
rect 8116 4496 8168 4548
rect 9496 4496 9548 4548
rect 11152 4564 11204 4616
rect 14280 4632 14332 4684
rect 15016 4632 15068 4684
rect 16028 4675 16080 4684
rect 16028 4641 16037 4675
rect 16037 4641 16071 4675
rect 16071 4641 16080 4675
rect 16028 4632 16080 4641
rect 17776 4675 17828 4684
rect 17776 4641 17785 4675
rect 17785 4641 17819 4675
rect 17819 4641 17828 4675
rect 17776 4632 17828 4641
rect 18144 4632 18196 4684
rect 18880 4632 18932 4684
rect 11428 4564 11480 4616
rect 11888 4564 11940 4616
rect 12072 4564 12124 4616
rect 13176 4564 13228 4616
rect 14372 4564 14424 4616
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 12716 4496 12768 4548
rect 13360 4496 13412 4548
rect 17132 4564 17184 4616
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 11152 4428 11204 4480
rect 12992 4428 13044 4480
rect 13636 4428 13688 4480
rect 15752 4428 15804 4480
rect 19064 4428 19116 4480
rect 20168 4428 20220 4480
rect 1782 4326 1834 4378
rect 1846 4326 1898 4378
rect 1910 4326 1962 4378
rect 1974 4326 2026 4378
rect 4782 4326 4834 4378
rect 4846 4326 4898 4378
rect 4910 4326 4962 4378
rect 4974 4326 5026 4378
rect 7782 4326 7834 4378
rect 7846 4326 7898 4378
rect 7910 4326 7962 4378
rect 7974 4326 8026 4378
rect 10782 4326 10834 4378
rect 10846 4326 10898 4378
rect 10910 4326 10962 4378
rect 10974 4326 11026 4378
rect 13782 4326 13834 4378
rect 13846 4326 13898 4378
rect 13910 4326 13962 4378
rect 13974 4326 14026 4378
rect 16782 4326 16834 4378
rect 16846 4326 16898 4378
rect 16910 4326 16962 4378
rect 16974 4326 17026 4378
rect 19782 4326 19834 4378
rect 19846 4326 19898 4378
rect 19910 4326 19962 4378
rect 19974 4326 20026 4378
rect 22782 4326 22834 4378
rect 22846 4326 22898 4378
rect 22910 4326 22962 4378
rect 22974 4326 23026 4378
rect 25782 4326 25834 4378
rect 25846 4326 25898 4378
rect 25910 4326 25962 4378
rect 25974 4326 26026 4378
rect 11888 4224 11940 4276
rect 13544 4224 13596 4276
rect 16028 4224 16080 4276
rect 16304 4224 16356 4276
rect 19616 4224 19668 4276
rect 6736 4156 6788 4208
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 8852 4156 8904 4208
rect 9036 4156 9088 4208
rect 10232 4156 10284 4208
rect 11796 4156 11848 4208
rect 12900 4156 12952 4208
rect 12992 4156 13044 4208
rect 16856 4156 16908 4208
rect 11152 4088 11204 4140
rect 8576 4063 8628 4072
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 6644 3884 6696 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 8300 3884 8352 3936
rect 9588 3884 9640 3936
rect 12716 4020 12768 4072
rect 14372 4088 14424 4140
rect 17500 4088 17552 4140
rect 17960 4088 18012 4140
rect 18604 4156 18656 4208
rect 18880 4088 18932 4140
rect 19616 4131 19668 4140
rect 19616 4097 19625 4131
rect 19625 4097 19659 4131
rect 19659 4097 19668 4131
rect 19616 4088 19668 4097
rect 14924 4020 14976 4072
rect 17776 4020 17828 4072
rect 13176 3952 13228 4004
rect 14464 3995 14516 4004
rect 14464 3961 14488 3995
rect 14488 3961 14516 3995
rect 16580 3995 16632 4004
rect 14464 3952 14516 3961
rect 16580 3961 16589 3995
rect 16589 3961 16623 3995
rect 16623 3961 16632 3995
rect 16580 3952 16632 3961
rect 17132 3952 17184 4004
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 19340 3952 19392 4004
rect 20444 3927 20496 3936
rect 20444 3893 20453 3927
rect 20453 3893 20487 3927
rect 20487 3893 20496 3927
rect 20444 3884 20496 3893
rect 3282 3782 3334 3834
rect 3346 3782 3398 3834
rect 3410 3782 3462 3834
rect 3474 3782 3526 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 6410 3782 6462 3834
rect 6474 3782 6526 3834
rect 9282 3782 9334 3834
rect 9346 3782 9398 3834
rect 9410 3782 9462 3834
rect 9474 3782 9526 3834
rect 12282 3782 12334 3834
rect 12346 3782 12398 3834
rect 12410 3782 12462 3834
rect 12474 3782 12526 3834
rect 15282 3782 15334 3834
rect 15346 3782 15398 3834
rect 15410 3782 15462 3834
rect 15474 3782 15526 3834
rect 18282 3782 18334 3834
rect 18346 3782 18398 3834
rect 18410 3782 18462 3834
rect 18474 3782 18526 3834
rect 21282 3782 21334 3834
rect 21346 3782 21398 3834
rect 21410 3782 21462 3834
rect 21474 3782 21526 3834
rect 24282 3782 24334 3834
rect 24346 3782 24398 3834
rect 24410 3782 24462 3834
rect 24474 3782 24526 3834
rect 27282 3782 27334 3834
rect 27346 3782 27398 3834
rect 27410 3782 27462 3834
rect 27474 3782 27526 3834
rect 7196 3680 7248 3732
rect 11428 3680 11480 3732
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 12900 3680 12952 3732
rect 14096 3680 14148 3732
rect 17960 3680 18012 3732
rect 19340 3680 19392 3732
rect 20168 3680 20220 3732
rect 8024 3612 8076 3664
rect 7656 3544 7708 3596
rect 8484 3544 8536 3596
rect 11336 3612 11388 3664
rect 14464 3612 14516 3664
rect 16856 3612 16908 3664
rect 8300 3476 8352 3528
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11428 3587 11480 3596
rect 11428 3553 11437 3587
rect 11437 3553 11471 3587
rect 11471 3553 11480 3587
rect 11428 3544 11480 3553
rect 14280 3544 14332 3596
rect 17500 3587 17552 3596
rect 17500 3553 17509 3587
rect 17509 3553 17543 3587
rect 17543 3553 17552 3587
rect 17500 3544 17552 3553
rect 8484 3408 8536 3460
rect 9772 3408 9824 3460
rect 12900 3476 12952 3528
rect 15752 3519 15804 3528
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 8852 3340 8904 3392
rect 9496 3340 9548 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 17132 3408 17184 3460
rect 14188 3340 14240 3392
rect 17960 3340 18012 3392
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 1782 3238 1834 3290
rect 1846 3238 1898 3290
rect 1910 3238 1962 3290
rect 1974 3238 2026 3290
rect 4782 3238 4834 3290
rect 4846 3238 4898 3290
rect 4910 3238 4962 3290
rect 4974 3238 5026 3290
rect 7782 3238 7834 3290
rect 7846 3238 7898 3290
rect 7910 3238 7962 3290
rect 7974 3238 8026 3290
rect 10782 3238 10834 3290
rect 10846 3238 10898 3290
rect 10910 3238 10962 3290
rect 10974 3238 11026 3290
rect 13782 3238 13834 3290
rect 13846 3238 13898 3290
rect 13910 3238 13962 3290
rect 13974 3238 14026 3290
rect 16782 3238 16834 3290
rect 16846 3238 16898 3290
rect 16910 3238 16962 3290
rect 16974 3238 17026 3290
rect 19782 3238 19834 3290
rect 19846 3238 19898 3290
rect 19910 3238 19962 3290
rect 19974 3238 20026 3290
rect 22782 3238 22834 3290
rect 22846 3238 22898 3290
rect 22910 3238 22962 3290
rect 22974 3238 23026 3290
rect 25782 3238 25834 3290
rect 25846 3238 25898 3290
rect 25910 3238 25962 3290
rect 25974 3238 26026 3290
rect 6644 3136 6696 3188
rect 8116 3136 8168 3188
rect 8576 3136 8628 3188
rect 9036 3136 9088 3188
rect 11428 3136 11480 3188
rect 9772 3111 9824 3120
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 10232 3068 10284 3120
rect 13084 3136 13136 3188
rect 16120 3136 16172 3188
rect 18604 3136 18656 3188
rect 20444 3136 20496 3188
rect 12624 3068 12676 3120
rect 13268 3068 13320 3120
rect 13636 3068 13688 3120
rect 14924 3111 14976 3120
rect 14924 3077 14933 3111
rect 14933 3077 14967 3111
rect 14967 3077 14976 3111
rect 14924 3068 14976 3077
rect 15016 3068 15068 3120
rect 18696 3111 18748 3120
rect 18696 3077 18705 3111
rect 18705 3077 18739 3111
rect 18739 3077 18748 3111
rect 18696 3068 18748 3077
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 7380 3000 7432 3052
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17960 3000 18012 3052
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 15752 2975 15804 2984
rect 12900 2932 12952 2941
rect 15752 2941 15761 2975
rect 15761 2941 15795 2975
rect 15795 2941 15804 2975
rect 15752 2932 15804 2941
rect 14372 2864 14424 2916
rect 13820 2796 13872 2848
rect 14188 2796 14240 2848
rect 17132 2796 17184 2848
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 3282 2694 3334 2746
rect 3346 2694 3398 2746
rect 3410 2694 3462 2746
rect 3474 2694 3526 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 6410 2694 6462 2746
rect 6474 2694 6526 2746
rect 9282 2694 9334 2746
rect 9346 2694 9398 2746
rect 9410 2694 9462 2746
rect 9474 2694 9526 2746
rect 12282 2694 12334 2746
rect 12346 2694 12398 2746
rect 12410 2694 12462 2746
rect 12474 2694 12526 2746
rect 15282 2694 15334 2746
rect 15346 2694 15398 2746
rect 15410 2694 15462 2746
rect 15474 2694 15526 2746
rect 18282 2694 18334 2746
rect 18346 2694 18398 2746
rect 18410 2694 18462 2746
rect 18474 2694 18526 2746
rect 21282 2694 21334 2746
rect 21346 2694 21398 2746
rect 21410 2694 21462 2746
rect 21474 2694 21526 2746
rect 24282 2694 24334 2746
rect 24346 2694 24398 2746
rect 24410 2694 24462 2746
rect 24474 2694 24526 2746
rect 27282 2694 27334 2746
rect 27346 2694 27398 2746
rect 27410 2694 27462 2746
rect 27474 2694 27526 2746
rect 7656 2635 7708 2644
rect 7656 2601 7665 2635
rect 7665 2601 7699 2635
rect 7699 2601 7708 2635
rect 7656 2592 7708 2601
rect 9772 2592 9824 2644
rect 10232 2592 10284 2644
rect 11244 2592 11296 2644
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 13268 2635 13320 2644
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 13360 2592 13412 2644
rect 13636 2524 13688 2576
rect 17500 2592 17552 2644
rect 14556 2524 14608 2576
rect 17960 2567 18012 2576
rect 17960 2533 17969 2567
rect 17969 2533 18003 2567
rect 18003 2533 18012 2567
rect 17960 2524 18012 2533
rect 7288 2388 7340 2440
rect 10048 2388 10100 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 14096 2431 14148 2440
rect 13820 2388 13872 2397
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 9128 2320 9180 2372
rect 16948 2320 17000 2372
rect 18236 2320 18288 2372
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9588 2252 9640 2304
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 1782 2150 1834 2202
rect 1846 2150 1898 2202
rect 1910 2150 1962 2202
rect 1974 2150 2026 2202
rect 4782 2150 4834 2202
rect 4846 2150 4898 2202
rect 4910 2150 4962 2202
rect 4974 2150 5026 2202
rect 7782 2150 7834 2202
rect 7846 2150 7898 2202
rect 7910 2150 7962 2202
rect 7974 2150 8026 2202
rect 10782 2150 10834 2202
rect 10846 2150 10898 2202
rect 10910 2150 10962 2202
rect 10974 2150 11026 2202
rect 13782 2150 13834 2202
rect 13846 2150 13898 2202
rect 13910 2150 13962 2202
rect 13974 2150 14026 2202
rect 16782 2150 16834 2202
rect 16846 2150 16898 2202
rect 16910 2150 16962 2202
rect 16974 2150 17026 2202
rect 19782 2150 19834 2202
rect 19846 2150 19898 2202
rect 19910 2150 19962 2202
rect 19974 2150 20026 2202
rect 22782 2150 22834 2202
rect 22846 2150 22898 2202
rect 22910 2150 22962 2202
rect 22974 2150 23026 2202
rect 25782 2150 25834 2202
rect 25846 2150 25898 2202
rect 25910 2150 25962 2202
rect 25974 2150 26026 2202
rect 20 8 72 60
rect 9956 8 10008 60
<< metal2 >>
rect 6366 30864 6422 31664
rect 15658 30864 15714 31664
rect 24858 30954 24914 31664
rect 24596 30926 24914 30954
rect 1756 29404 2052 29424
rect 1812 29402 1836 29404
rect 1892 29402 1916 29404
rect 1972 29402 1996 29404
rect 1834 29350 1836 29402
rect 1898 29350 1910 29402
rect 1972 29350 1974 29402
rect 1812 29348 1836 29350
rect 1892 29348 1916 29350
rect 1972 29348 1996 29350
rect 1756 29328 2052 29348
rect 4756 29404 5052 29424
rect 4812 29402 4836 29404
rect 4892 29402 4916 29404
rect 4972 29402 4996 29404
rect 4834 29350 4836 29402
rect 4898 29350 4910 29402
rect 4972 29350 4974 29402
rect 4812 29348 4836 29350
rect 4892 29348 4916 29350
rect 4972 29348 4996 29350
rect 4756 29328 5052 29348
rect 7756 29404 8052 29424
rect 7812 29402 7836 29404
rect 7892 29402 7916 29404
rect 7972 29402 7996 29404
rect 7834 29350 7836 29402
rect 7898 29350 7910 29402
rect 7972 29350 7974 29402
rect 7812 29348 7836 29350
rect 7892 29348 7916 29350
rect 7972 29348 7996 29350
rect 7756 29328 8052 29348
rect 10756 29404 11052 29424
rect 10812 29402 10836 29404
rect 10892 29402 10916 29404
rect 10972 29402 10996 29404
rect 10834 29350 10836 29402
rect 10898 29350 10910 29402
rect 10972 29350 10974 29402
rect 10812 29348 10836 29350
rect 10892 29348 10916 29350
rect 10972 29348 10996 29350
rect 10756 29328 11052 29348
rect 13756 29404 14052 29424
rect 13812 29402 13836 29404
rect 13892 29402 13916 29404
rect 13972 29402 13996 29404
rect 13834 29350 13836 29402
rect 13898 29350 13910 29402
rect 13972 29350 13974 29402
rect 13812 29348 13836 29350
rect 13892 29348 13916 29350
rect 13972 29348 13996 29350
rect 13756 29328 14052 29348
rect 16756 29404 17052 29424
rect 16812 29402 16836 29404
rect 16892 29402 16916 29404
rect 16972 29402 16996 29404
rect 16834 29350 16836 29402
rect 16898 29350 16910 29402
rect 16972 29350 16974 29402
rect 16812 29348 16836 29350
rect 16892 29348 16916 29350
rect 16972 29348 16996 29350
rect 16756 29328 17052 29348
rect 19756 29404 20052 29424
rect 19812 29402 19836 29404
rect 19892 29402 19916 29404
rect 19972 29402 19996 29404
rect 19834 29350 19836 29402
rect 19898 29350 19910 29402
rect 19972 29350 19974 29402
rect 19812 29348 19836 29350
rect 19892 29348 19916 29350
rect 19972 29348 19996 29350
rect 19756 29328 20052 29348
rect 22756 29404 23052 29424
rect 22812 29402 22836 29404
rect 22892 29402 22916 29404
rect 22972 29402 22996 29404
rect 22834 29350 22836 29402
rect 22898 29350 22910 29402
rect 22972 29350 22974 29402
rect 22812 29348 22836 29350
rect 22892 29348 22916 29350
rect 22972 29348 22996 29350
rect 22756 29328 23052 29348
rect 3256 28860 3552 28880
rect 3312 28858 3336 28860
rect 3392 28858 3416 28860
rect 3472 28858 3496 28860
rect 3334 28806 3336 28858
rect 3398 28806 3410 28858
rect 3472 28806 3474 28858
rect 3312 28804 3336 28806
rect 3392 28804 3416 28806
rect 3472 28804 3496 28806
rect 3256 28784 3552 28804
rect 6256 28860 6552 28880
rect 6312 28858 6336 28860
rect 6392 28858 6416 28860
rect 6472 28858 6496 28860
rect 6334 28806 6336 28858
rect 6398 28806 6410 28858
rect 6472 28806 6474 28858
rect 6312 28804 6336 28806
rect 6392 28804 6416 28806
rect 6472 28804 6496 28806
rect 6256 28784 6552 28804
rect 9256 28860 9552 28880
rect 9312 28858 9336 28860
rect 9392 28858 9416 28860
rect 9472 28858 9496 28860
rect 9334 28806 9336 28858
rect 9398 28806 9410 28858
rect 9472 28806 9474 28858
rect 9312 28804 9336 28806
rect 9392 28804 9416 28806
rect 9472 28804 9496 28806
rect 9256 28784 9552 28804
rect 12256 28860 12552 28880
rect 12312 28858 12336 28860
rect 12392 28858 12416 28860
rect 12472 28858 12496 28860
rect 12334 28806 12336 28858
rect 12398 28806 12410 28858
rect 12472 28806 12474 28858
rect 12312 28804 12336 28806
rect 12392 28804 12416 28806
rect 12472 28804 12496 28806
rect 12256 28784 12552 28804
rect 15256 28860 15552 28880
rect 15312 28858 15336 28860
rect 15392 28858 15416 28860
rect 15472 28858 15496 28860
rect 15334 28806 15336 28858
rect 15398 28806 15410 28858
rect 15472 28806 15474 28858
rect 15312 28804 15336 28806
rect 15392 28804 15416 28806
rect 15472 28804 15496 28806
rect 15256 28784 15552 28804
rect 18256 28860 18552 28880
rect 18312 28858 18336 28860
rect 18392 28858 18416 28860
rect 18472 28858 18496 28860
rect 18334 28806 18336 28858
rect 18398 28806 18410 28858
rect 18472 28806 18474 28858
rect 18312 28804 18336 28806
rect 18392 28804 18416 28806
rect 18472 28804 18496 28806
rect 18256 28784 18552 28804
rect 21256 28860 21552 28880
rect 21312 28858 21336 28860
rect 21392 28858 21416 28860
rect 21472 28858 21496 28860
rect 21334 28806 21336 28858
rect 21398 28806 21410 28858
rect 21472 28806 21474 28858
rect 21312 28804 21336 28806
rect 21392 28804 21416 28806
rect 21472 28804 21496 28806
rect 21256 28784 21552 28804
rect 24256 28860 24552 28880
rect 24312 28858 24336 28860
rect 24392 28858 24416 28860
rect 24472 28858 24496 28860
rect 24334 28806 24336 28858
rect 24398 28806 24410 28858
rect 24472 28806 24474 28858
rect 24312 28804 24336 28806
rect 24392 28804 24416 28806
rect 24472 28804 24496 28806
rect 24256 28784 24552 28804
rect 1756 28316 2052 28336
rect 1812 28314 1836 28316
rect 1892 28314 1916 28316
rect 1972 28314 1996 28316
rect 1834 28262 1836 28314
rect 1898 28262 1910 28314
rect 1972 28262 1974 28314
rect 1812 28260 1836 28262
rect 1892 28260 1916 28262
rect 1972 28260 1996 28262
rect 1756 28240 2052 28260
rect 4756 28316 5052 28336
rect 4812 28314 4836 28316
rect 4892 28314 4916 28316
rect 4972 28314 4996 28316
rect 4834 28262 4836 28314
rect 4898 28262 4910 28314
rect 4972 28262 4974 28314
rect 4812 28260 4836 28262
rect 4892 28260 4916 28262
rect 4972 28260 4996 28262
rect 4756 28240 5052 28260
rect 7756 28316 8052 28336
rect 7812 28314 7836 28316
rect 7892 28314 7916 28316
rect 7972 28314 7996 28316
rect 7834 28262 7836 28314
rect 7898 28262 7910 28314
rect 7972 28262 7974 28314
rect 7812 28260 7836 28262
rect 7892 28260 7916 28262
rect 7972 28260 7996 28262
rect 7756 28240 8052 28260
rect 10756 28316 11052 28336
rect 10812 28314 10836 28316
rect 10892 28314 10916 28316
rect 10972 28314 10996 28316
rect 10834 28262 10836 28314
rect 10898 28262 10910 28314
rect 10972 28262 10974 28314
rect 10812 28260 10836 28262
rect 10892 28260 10916 28262
rect 10972 28260 10996 28262
rect 10756 28240 11052 28260
rect 13756 28316 14052 28336
rect 13812 28314 13836 28316
rect 13892 28314 13916 28316
rect 13972 28314 13996 28316
rect 13834 28262 13836 28314
rect 13898 28262 13910 28314
rect 13972 28262 13974 28314
rect 13812 28260 13836 28262
rect 13892 28260 13916 28262
rect 13972 28260 13996 28262
rect 13756 28240 14052 28260
rect 16756 28316 17052 28336
rect 16812 28314 16836 28316
rect 16892 28314 16916 28316
rect 16972 28314 16996 28316
rect 16834 28262 16836 28314
rect 16898 28262 16910 28314
rect 16972 28262 16974 28314
rect 16812 28260 16836 28262
rect 16892 28260 16916 28262
rect 16972 28260 16996 28262
rect 16756 28240 17052 28260
rect 19756 28316 20052 28336
rect 19812 28314 19836 28316
rect 19892 28314 19916 28316
rect 19972 28314 19996 28316
rect 19834 28262 19836 28314
rect 19898 28262 19910 28314
rect 19972 28262 19974 28314
rect 19812 28260 19836 28262
rect 19892 28260 19916 28262
rect 19972 28260 19996 28262
rect 19756 28240 20052 28260
rect 22756 28316 23052 28336
rect 22812 28314 22836 28316
rect 22892 28314 22916 28316
rect 22972 28314 22996 28316
rect 22834 28262 22836 28314
rect 22898 28262 22910 28314
rect 22972 28262 22974 28314
rect 22812 28260 22836 28262
rect 22892 28260 22916 28262
rect 22972 28260 22996 28262
rect 22756 28240 23052 28260
rect 3256 27772 3552 27792
rect 3312 27770 3336 27772
rect 3392 27770 3416 27772
rect 3472 27770 3496 27772
rect 3334 27718 3336 27770
rect 3398 27718 3410 27770
rect 3472 27718 3474 27770
rect 3312 27716 3336 27718
rect 3392 27716 3416 27718
rect 3472 27716 3496 27718
rect 3256 27696 3552 27716
rect 6256 27772 6552 27792
rect 6312 27770 6336 27772
rect 6392 27770 6416 27772
rect 6472 27770 6496 27772
rect 6334 27718 6336 27770
rect 6398 27718 6410 27770
rect 6472 27718 6474 27770
rect 6312 27716 6336 27718
rect 6392 27716 6416 27718
rect 6472 27716 6496 27718
rect 6256 27696 6552 27716
rect 9256 27772 9552 27792
rect 9312 27770 9336 27772
rect 9392 27770 9416 27772
rect 9472 27770 9496 27772
rect 9334 27718 9336 27770
rect 9398 27718 9410 27770
rect 9472 27718 9474 27770
rect 9312 27716 9336 27718
rect 9392 27716 9416 27718
rect 9472 27716 9496 27718
rect 9256 27696 9552 27716
rect 12256 27772 12552 27792
rect 12312 27770 12336 27772
rect 12392 27770 12416 27772
rect 12472 27770 12496 27772
rect 12334 27718 12336 27770
rect 12398 27718 12410 27770
rect 12472 27718 12474 27770
rect 12312 27716 12336 27718
rect 12392 27716 12416 27718
rect 12472 27716 12496 27718
rect 12256 27696 12552 27716
rect 15256 27772 15552 27792
rect 15312 27770 15336 27772
rect 15392 27770 15416 27772
rect 15472 27770 15496 27772
rect 15334 27718 15336 27770
rect 15398 27718 15410 27770
rect 15472 27718 15474 27770
rect 15312 27716 15336 27718
rect 15392 27716 15416 27718
rect 15472 27716 15496 27718
rect 15256 27696 15552 27716
rect 18256 27772 18552 27792
rect 18312 27770 18336 27772
rect 18392 27770 18416 27772
rect 18472 27770 18496 27772
rect 18334 27718 18336 27770
rect 18398 27718 18410 27770
rect 18472 27718 18474 27770
rect 18312 27716 18336 27718
rect 18392 27716 18416 27718
rect 18472 27716 18496 27718
rect 18256 27696 18552 27716
rect 21256 27772 21552 27792
rect 21312 27770 21336 27772
rect 21392 27770 21416 27772
rect 21472 27770 21496 27772
rect 21334 27718 21336 27770
rect 21398 27718 21410 27770
rect 21472 27718 21474 27770
rect 21312 27716 21336 27718
rect 21392 27716 21416 27718
rect 21472 27716 21496 27718
rect 21256 27696 21552 27716
rect 24256 27772 24552 27792
rect 24312 27770 24336 27772
rect 24392 27770 24416 27772
rect 24472 27770 24496 27772
rect 24334 27718 24336 27770
rect 24398 27718 24410 27770
rect 24472 27718 24474 27770
rect 24312 27716 24336 27718
rect 24392 27716 24416 27718
rect 24472 27716 24496 27718
rect 24256 27696 24552 27716
rect 24596 27470 24624 30926
rect 24858 30864 24914 30926
rect 25756 29404 26052 29424
rect 25812 29402 25836 29404
rect 25892 29402 25916 29404
rect 25972 29402 25996 29404
rect 25834 29350 25836 29402
rect 25898 29350 25910 29402
rect 25972 29350 25974 29402
rect 25812 29348 25836 29350
rect 25892 29348 25916 29350
rect 25972 29348 25996 29350
rect 25756 29328 26052 29348
rect 27256 28860 27552 28880
rect 27312 28858 27336 28860
rect 27392 28858 27416 28860
rect 27472 28858 27496 28860
rect 27334 28806 27336 28858
rect 27398 28806 27410 28858
rect 27472 28806 27474 28858
rect 27312 28804 27336 28806
rect 27392 28804 27416 28806
rect 27472 28804 27496 28806
rect 27256 28784 27552 28804
rect 25756 28316 26052 28336
rect 25812 28314 25836 28316
rect 25892 28314 25916 28316
rect 25972 28314 25996 28316
rect 25834 28262 25836 28314
rect 25898 28262 25910 28314
rect 25972 28262 25974 28314
rect 25812 28260 25836 28262
rect 25892 28260 25916 28262
rect 25972 28260 25996 28262
rect 25756 28240 26052 28260
rect 27256 27772 27552 27792
rect 27312 27770 27336 27772
rect 27392 27770 27416 27772
rect 27472 27770 27496 27772
rect 27334 27718 27336 27770
rect 27398 27718 27410 27770
rect 27472 27718 27474 27770
rect 27312 27716 27336 27718
rect 27392 27716 27416 27718
rect 27472 27716 27496 27718
rect 27256 27696 27552 27716
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 21640 27396 21692 27402
rect 21640 27338 21692 27344
rect 1756 27228 2052 27248
rect 1812 27226 1836 27228
rect 1892 27226 1916 27228
rect 1972 27226 1996 27228
rect 1834 27174 1836 27226
rect 1898 27174 1910 27226
rect 1972 27174 1974 27226
rect 1812 27172 1836 27174
rect 1892 27172 1916 27174
rect 1972 27172 1996 27174
rect 1756 27152 2052 27172
rect 4756 27228 5052 27248
rect 4812 27226 4836 27228
rect 4892 27226 4916 27228
rect 4972 27226 4996 27228
rect 4834 27174 4836 27226
rect 4898 27174 4910 27226
rect 4972 27174 4974 27226
rect 4812 27172 4836 27174
rect 4892 27172 4916 27174
rect 4972 27172 4996 27174
rect 4756 27152 5052 27172
rect 7756 27228 8052 27248
rect 7812 27226 7836 27228
rect 7892 27226 7916 27228
rect 7972 27226 7996 27228
rect 7834 27174 7836 27226
rect 7898 27174 7910 27226
rect 7972 27174 7974 27226
rect 7812 27172 7836 27174
rect 7892 27172 7916 27174
rect 7972 27172 7996 27174
rect 7756 27152 8052 27172
rect 10756 27228 11052 27248
rect 10812 27226 10836 27228
rect 10892 27226 10916 27228
rect 10972 27226 10996 27228
rect 10834 27174 10836 27226
rect 10898 27174 10910 27226
rect 10972 27174 10974 27226
rect 10812 27172 10836 27174
rect 10892 27172 10916 27174
rect 10972 27172 10996 27174
rect 10756 27152 11052 27172
rect 13756 27228 14052 27248
rect 13812 27226 13836 27228
rect 13892 27226 13916 27228
rect 13972 27226 13996 27228
rect 13834 27174 13836 27226
rect 13898 27174 13910 27226
rect 13972 27174 13974 27226
rect 13812 27172 13836 27174
rect 13892 27172 13916 27174
rect 13972 27172 13996 27174
rect 13756 27152 14052 27172
rect 16756 27228 17052 27248
rect 16812 27226 16836 27228
rect 16892 27226 16916 27228
rect 16972 27226 16996 27228
rect 16834 27174 16836 27226
rect 16898 27174 16910 27226
rect 16972 27174 16974 27226
rect 16812 27172 16836 27174
rect 16892 27172 16916 27174
rect 16972 27172 16996 27174
rect 16756 27152 17052 27172
rect 19756 27228 20052 27248
rect 19812 27226 19836 27228
rect 19892 27226 19916 27228
rect 19972 27226 19996 27228
rect 19834 27174 19836 27226
rect 19898 27174 19910 27226
rect 19972 27174 19974 27226
rect 19812 27172 19836 27174
rect 19892 27172 19916 27174
rect 19972 27172 19996 27174
rect 19756 27152 20052 27172
rect 3256 26684 3552 26704
rect 3312 26682 3336 26684
rect 3392 26682 3416 26684
rect 3472 26682 3496 26684
rect 3334 26630 3336 26682
rect 3398 26630 3410 26682
rect 3472 26630 3474 26682
rect 3312 26628 3336 26630
rect 3392 26628 3416 26630
rect 3472 26628 3496 26630
rect 3256 26608 3552 26628
rect 6256 26684 6552 26704
rect 6312 26682 6336 26684
rect 6392 26682 6416 26684
rect 6472 26682 6496 26684
rect 6334 26630 6336 26682
rect 6398 26630 6410 26682
rect 6472 26630 6474 26682
rect 6312 26628 6336 26630
rect 6392 26628 6416 26630
rect 6472 26628 6496 26630
rect 6256 26608 6552 26628
rect 9256 26684 9552 26704
rect 9312 26682 9336 26684
rect 9392 26682 9416 26684
rect 9472 26682 9496 26684
rect 9334 26630 9336 26682
rect 9398 26630 9410 26682
rect 9472 26630 9474 26682
rect 9312 26628 9336 26630
rect 9392 26628 9416 26630
rect 9472 26628 9496 26630
rect 9256 26608 9552 26628
rect 12256 26684 12552 26704
rect 12312 26682 12336 26684
rect 12392 26682 12416 26684
rect 12472 26682 12496 26684
rect 12334 26630 12336 26682
rect 12398 26630 12410 26682
rect 12472 26630 12474 26682
rect 12312 26628 12336 26630
rect 12392 26628 12416 26630
rect 12472 26628 12496 26630
rect 12256 26608 12552 26628
rect 15256 26684 15552 26704
rect 15312 26682 15336 26684
rect 15392 26682 15416 26684
rect 15472 26682 15496 26684
rect 15334 26630 15336 26682
rect 15398 26630 15410 26682
rect 15472 26630 15474 26682
rect 15312 26628 15336 26630
rect 15392 26628 15416 26630
rect 15472 26628 15496 26630
rect 15256 26608 15552 26628
rect 18256 26684 18552 26704
rect 18312 26682 18336 26684
rect 18392 26682 18416 26684
rect 18472 26682 18496 26684
rect 18334 26630 18336 26682
rect 18398 26630 18410 26682
rect 18472 26630 18474 26682
rect 18312 26628 18336 26630
rect 18392 26628 18416 26630
rect 18472 26628 18496 26630
rect 18256 26608 18552 26628
rect 21256 26684 21552 26704
rect 21312 26682 21336 26684
rect 21392 26682 21416 26684
rect 21472 26682 21496 26684
rect 21334 26630 21336 26682
rect 21398 26630 21410 26682
rect 21472 26630 21474 26682
rect 21312 26628 21336 26630
rect 21392 26628 21416 26630
rect 21472 26628 21496 26630
rect 21256 26608 21552 26628
rect 1756 26140 2052 26160
rect 1812 26138 1836 26140
rect 1892 26138 1916 26140
rect 1972 26138 1996 26140
rect 1834 26086 1836 26138
rect 1898 26086 1910 26138
rect 1972 26086 1974 26138
rect 1812 26084 1836 26086
rect 1892 26084 1916 26086
rect 1972 26084 1996 26086
rect 1756 26064 2052 26084
rect 4756 26140 5052 26160
rect 4812 26138 4836 26140
rect 4892 26138 4916 26140
rect 4972 26138 4996 26140
rect 4834 26086 4836 26138
rect 4898 26086 4910 26138
rect 4972 26086 4974 26138
rect 4812 26084 4836 26086
rect 4892 26084 4916 26086
rect 4972 26084 4996 26086
rect 4756 26064 5052 26084
rect 7756 26140 8052 26160
rect 7812 26138 7836 26140
rect 7892 26138 7916 26140
rect 7972 26138 7996 26140
rect 7834 26086 7836 26138
rect 7898 26086 7910 26138
rect 7972 26086 7974 26138
rect 7812 26084 7836 26086
rect 7892 26084 7916 26086
rect 7972 26084 7996 26086
rect 7756 26064 8052 26084
rect 10756 26140 11052 26160
rect 10812 26138 10836 26140
rect 10892 26138 10916 26140
rect 10972 26138 10996 26140
rect 10834 26086 10836 26138
rect 10898 26086 10910 26138
rect 10972 26086 10974 26138
rect 10812 26084 10836 26086
rect 10892 26084 10916 26086
rect 10972 26084 10996 26086
rect 10756 26064 11052 26084
rect 13756 26140 14052 26160
rect 13812 26138 13836 26140
rect 13892 26138 13916 26140
rect 13972 26138 13996 26140
rect 13834 26086 13836 26138
rect 13898 26086 13910 26138
rect 13972 26086 13974 26138
rect 13812 26084 13836 26086
rect 13892 26084 13916 26086
rect 13972 26084 13996 26086
rect 13756 26064 14052 26084
rect 16756 26140 17052 26160
rect 16812 26138 16836 26140
rect 16892 26138 16916 26140
rect 16972 26138 16996 26140
rect 16834 26086 16836 26138
rect 16898 26086 16910 26138
rect 16972 26086 16974 26138
rect 16812 26084 16836 26086
rect 16892 26084 16916 26086
rect 16972 26084 16996 26086
rect 16756 26064 17052 26084
rect 19756 26140 20052 26160
rect 19812 26138 19836 26140
rect 19892 26138 19916 26140
rect 19972 26138 19996 26140
rect 19834 26086 19836 26138
rect 19898 26086 19910 26138
rect 19972 26086 19974 26138
rect 19812 26084 19836 26086
rect 19892 26084 19916 26086
rect 19972 26084 19996 26086
rect 19756 26064 20052 26084
rect 3256 25596 3552 25616
rect 3312 25594 3336 25596
rect 3392 25594 3416 25596
rect 3472 25594 3496 25596
rect 3334 25542 3336 25594
rect 3398 25542 3410 25594
rect 3472 25542 3474 25594
rect 3312 25540 3336 25542
rect 3392 25540 3416 25542
rect 3472 25540 3496 25542
rect 3256 25520 3552 25540
rect 6256 25596 6552 25616
rect 6312 25594 6336 25596
rect 6392 25594 6416 25596
rect 6472 25594 6496 25596
rect 6334 25542 6336 25594
rect 6398 25542 6410 25594
rect 6472 25542 6474 25594
rect 6312 25540 6336 25542
rect 6392 25540 6416 25542
rect 6472 25540 6496 25542
rect 6256 25520 6552 25540
rect 9256 25596 9552 25616
rect 9312 25594 9336 25596
rect 9392 25594 9416 25596
rect 9472 25594 9496 25596
rect 9334 25542 9336 25594
rect 9398 25542 9410 25594
rect 9472 25542 9474 25594
rect 9312 25540 9336 25542
rect 9392 25540 9416 25542
rect 9472 25540 9496 25542
rect 9256 25520 9552 25540
rect 12256 25596 12552 25616
rect 12312 25594 12336 25596
rect 12392 25594 12416 25596
rect 12472 25594 12496 25596
rect 12334 25542 12336 25594
rect 12398 25542 12410 25594
rect 12472 25542 12474 25594
rect 12312 25540 12336 25542
rect 12392 25540 12416 25542
rect 12472 25540 12496 25542
rect 12256 25520 12552 25540
rect 15256 25596 15552 25616
rect 15312 25594 15336 25596
rect 15392 25594 15416 25596
rect 15472 25594 15496 25596
rect 15334 25542 15336 25594
rect 15398 25542 15410 25594
rect 15472 25542 15474 25594
rect 15312 25540 15336 25542
rect 15392 25540 15416 25542
rect 15472 25540 15496 25542
rect 15256 25520 15552 25540
rect 18256 25596 18552 25616
rect 18312 25594 18336 25596
rect 18392 25594 18416 25596
rect 18472 25594 18496 25596
rect 18334 25542 18336 25594
rect 18398 25542 18410 25594
rect 18472 25542 18474 25594
rect 18312 25540 18336 25542
rect 18392 25540 18416 25542
rect 18472 25540 18496 25542
rect 18256 25520 18552 25540
rect 21256 25596 21552 25616
rect 21312 25594 21336 25596
rect 21392 25594 21416 25596
rect 21472 25594 21496 25596
rect 21334 25542 21336 25594
rect 21398 25542 21410 25594
rect 21472 25542 21474 25594
rect 21312 25540 21336 25542
rect 21392 25540 21416 25542
rect 21472 25540 21496 25542
rect 21256 25520 21552 25540
rect 1756 25052 2052 25072
rect 1812 25050 1836 25052
rect 1892 25050 1916 25052
rect 1972 25050 1996 25052
rect 1834 24998 1836 25050
rect 1898 24998 1910 25050
rect 1972 24998 1974 25050
rect 1812 24996 1836 24998
rect 1892 24996 1916 24998
rect 1972 24996 1996 24998
rect 1756 24976 2052 24996
rect 4756 25052 5052 25072
rect 4812 25050 4836 25052
rect 4892 25050 4916 25052
rect 4972 25050 4996 25052
rect 4834 24998 4836 25050
rect 4898 24998 4910 25050
rect 4972 24998 4974 25050
rect 4812 24996 4836 24998
rect 4892 24996 4916 24998
rect 4972 24996 4996 24998
rect 4756 24976 5052 24996
rect 7756 25052 8052 25072
rect 7812 25050 7836 25052
rect 7892 25050 7916 25052
rect 7972 25050 7996 25052
rect 7834 24998 7836 25050
rect 7898 24998 7910 25050
rect 7972 24998 7974 25050
rect 7812 24996 7836 24998
rect 7892 24996 7916 24998
rect 7972 24996 7996 24998
rect 7756 24976 8052 24996
rect 10756 25052 11052 25072
rect 10812 25050 10836 25052
rect 10892 25050 10916 25052
rect 10972 25050 10996 25052
rect 10834 24998 10836 25050
rect 10898 24998 10910 25050
rect 10972 24998 10974 25050
rect 10812 24996 10836 24998
rect 10892 24996 10916 24998
rect 10972 24996 10996 24998
rect 10756 24976 11052 24996
rect 13756 25052 14052 25072
rect 13812 25050 13836 25052
rect 13892 25050 13916 25052
rect 13972 25050 13996 25052
rect 13834 24998 13836 25050
rect 13898 24998 13910 25050
rect 13972 24998 13974 25050
rect 13812 24996 13836 24998
rect 13892 24996 13916 24998
rect 13972 24996 13996 24998
rect 13756 24976 14052 24996
rect 16756 25052 17052 25072
rect 16812 25050 16836 25052
rect 16892 25050 16916 25052
rect 16972 25050 16996 25052
rect 16834 24998 16836 25050
rect 16898 24998 16910 25050
rect 16972 24998 16974 25050
rect 16812 24996 16836 24998
rect 16892 24996 16916 24998
rect 16972 24996 16996 24998
rect 16756 24976 17052 24996
rect 19756 25052 20052 25072
rect 19812 25050 19836 25052
rect 19892 25050 19916 25052
rect 19972 25050 19996 25052
rect 19834 24998 19836 25050
rect 19898 24998 19910 25050
rect 19972 24998 19974 25050
rect 19812 24996 19836 24998
rect 19892 24996 19916 24998
rect 19972 24996 19996 24998
rect 19756 24976 20052 24996
rect 3256 24508 3552 24528
rect 3312 24506 3336 24508
rect 3392 24506 3416 24508
rect 3472 24506 3496 24508
rect 3334 24454 3336 24506
rect 3398 24454 3410 24506
rect 3472 24454 3474 24506
rect 3312 24452 3336 24454
rect 3392 24452 3416 24454
rect 3472 24452 3496 24454
rect 3256 24432 3552 24452
rect 6256 24508 6552 24528
rect 6312 24506 6336 24508
rect 6392 24506 6416 24508
rect 6472 24506 6496 24508
rect 6334 24454 6336 24506
rect 6398 24454 6410 24506
rect 6472 24454 6474 24506
rect 6312 24452 6336 24454
rect 6392 24452 6416 24454
rect 6472 24452 6496 24454
rect 6256 24432 6552 24452
rect 9256 24508 9552 24528
rect 9312 24506 9336 24508
rect 9392 24506 9416 24508
rect 9472 24506 9496 24508
rect 9334 24454 9336 24506
rect 9398 24454 9410 24506
rect 9472 24454 9474 24506
rect 9312 24452 9336 24454
rect 9392 24452 9416 24454
rect 9472 24452 9496 24454
rect 9256 24432 9552 24452
rect 12256 24508 12552 24528
rect 12312 24506 12336 24508
rect 12392 24506 12416 24508
rect 12472 24506 12496 24508
rect 12334 24454 12336 24506
rect 12398 24454 12410 24506
rect 12472 24454 12474 24506
rect 12312 24452 12336 24454
rect 12392 24452 12416 24454
rect 12472 24452 12496 24454
rect 12256 24432 12552 24452
rect 15256 24508 15552 24528
rect 15312 24506 15336 24508
rect 15392 24506 15416 24508
rect 15472 24506 15496 24508
rect 15334 24454 15336 24506
rect 15398 24454 15410 24506
rect 15472 24454 15474 24506
rect 15312 24452 15336 24454
rect 15392 24452 15416 24454
rect 15472 24452 15496 24454
rect 15256 24432 15552 24452
rect 18256 24508 18552 24528
rect 18312 24506 18336 24508
rect 18392 24506 18416 24508
rect 18472 24506 18496 24508
rect 18334 24454 18336 24506
rect 18398 24454 18410 24506
rect 18472 24454 18474 24506
rect 18312 24452 18336 24454
rect 18392 24452 18416 24454
rect 18472 24452 18496 24454
rect 18256 24432 18552 24452
rect 21256 24508 21552 24528
rect 21312 24506 21336 24508
rect 21392 24506 21416 24508
rect 21472 24506 21496 24508
rect 21334 24454 21336 24506
rect 21398 24454 21410 24506
rect 21472 24454 21474 24506
rect 21312 24452 21336 24454
rect 21392 24452 21416 24454
rect 21472 24452 21496 24454
rect 21256 24432 21552 24452
rect 1756 23964 2052 23984
rect 1812 23962 1836 23964
rect 1892 23962 1916 23964
rect 1972 23962 1996 23964
rect 1834 23910 1836 23962
rect 1898 23910 1910 23962
rect 1972 23910 1974 23962
rect 1812 23908 1836 23910
rect 1892 23908 1916 23910
rect 1972 23908 1996 23910
rect 1756 23888 2052 23908
rect 4756 23964 5052 23984
rect 4812 23962 4836 23964
rect 4892 23962 4916 23964
rect 4972 23962 4996 23964
rect 4834 23910 4836 23962
rect 4898 23910 4910 23962
rect 4972 23910 4974 23962
rect 4812 23908 4836 23910
rect 4892 23908 4916 23910
rect 4972 23908 4996 23910
rect 4756 23888 5052 23908
rect 7756 23964 8052 23984
rect 7812 23962 7836 23964
rect 7892 23962 7916 23964
rect 7972 23962 7996 23964
rect 7834 23910 7836 23962
rect 7898 23910 7910 23962
rect 7972 23910 7974 23962
rect 7812 23908 7836 23910
rect 7892 23908 7916 23910
rect 7972 23908 7996 23910
rect 7756 23888 8052 23908
rect 10756 23964 11052 23984
rect 10812 23962 10836 23964
rect 10892 23962 10916 23964
rect 10972 23962 10996 23964
rect 10834 23910 10836 23962
rect 10898 23910 10910 23962
rect 10972 23910 10974 23962
rect 10812 23908 10836 23910
rect 10892 23908 10916 23910
rect 10972 23908 10996 23910
rect 10756 23888 11052 23908
rect 13756 23964 14052 23984
rect 13812 23962 13836 23964
rect 13892 23962 13916 23964
rect 13972 23962 13996 23964
rect 13834 23910 13836 23962
rect 13898 23910 13910 23962
rect 13972 23910 13974 23962
rect 13812 23908 13836 23910
rect 13892 23908 13916 23910
rect 13972 23908 13996 23910
rect 13756 23888 14052 23908
rect 16756 23964 17052 23984
rect 16812 23962 16836 23964
rect 16892 23962 16916 23964
rect 16972 23962 16996 23964
rect 16834 23910 16836 23962
rect 16898 23910 16910 23962
rect 16972 23910 16974 23962
rect 16812 23908 16836 23910
rect 16892 23908 16916 23910
rect 16972 23908 16996 23910
rect 16756 23888 17052 23908
rect 19756 23964 20052 23984
rect 19812 23962 19836 23964
rect 19892 23962 19916 23964
rect 19972 23962 19996 23964
rect 19834 23910 19836 23962
rect 19898 23910 19910 23962
rect 19972 23910 19974 23962
rect 19812 23908 19836 23910
rect 19892 23908 19916 23910
rect 19972 23908 19996 23910
rect 19756 23888 20052 23908
rect 3256 23420 3552 23440
rect 3312 23418 3336 23420
rect 3392 23418 3416 23420
rect 3472 23418 3496 23420
rect 3334 23366 3336 23418
rect 3398 23366 3410 23418
rect 3472 23366 3474 23418
rect 3312 23364 3336 23366
rect 3392 23364 3416 23366
rect 3472 23364 3496 23366
rect 3256 23344 3552 23364
rect 6256 23420 6552 23440
rect 6312 23418 6336 23420
rect 6392 23418 6416 23420
rect 6472 23418 6496 23420
rect 6334 23366 6336 23418
rect 6398 23366 6410 23418
rect 6472 23366 6474 23418
rect 6312 23364 6336 23366
rect 6392 23364 6416 23366
rect 6472 23364 6496 23366
rect 6256 23344 6552 23364
rect 9256 23420 9552 23440
rect 9312 23418 9336 23420
rect 9392 23418 9416 23420
rect 9472 23418 9496 23420
rect 9334 23366 9336 23418
rect 9398 23366 9410 23418
rect 9472 23366 9474 23418
rect 9312 23364 9336 23366
rect 9392 23364 9416 23366
rect 9472 23364 9496 23366
rect 9256 23344 9552 23364
rect 12256 23420 12552 23440
rect 12312 23418 12336 23420
rect 12392 23418 12416 23420
rect 12472 23418 12496 23420
rect 12334 23366 12336 23418
rect 12398 23366 12410 23418
rect 12472 23366 12474 23418
rect 12312 23364 12336 23366
rect 12392 23364 12416 23366
rect 12472 23364 12496 23366
rect 12256 23344 12552 23364
rect 15256 23420 15552 23440
rect 15312 23418 15336 23420
rect 15392 23418 15416 23420
rect 15472 23418 15496 23420
rect 15334 23366 15336 23418
rect 15398 23366 15410 23418
rect 15472 23366 15474 23418
rect 15312 23364 15336 23366
rect 15392 23364 15416 23366
rect 15472 23364 15496 23366
rect 15256 23344 15552 23364
rect 18256 23420 18552 23440
rect 18312 23418 18336 23420
rect 18392 23418 18416 23420
rect 18472 23418 18496 23420
rect 18334 23366 18336 23418
rect 18398 23366 18410 23418
rect 18472 23366 18474 23418
rect 18312 23364 18336 23366
rect 18392 23364 18416 23366
rect 18472 23364 18496 23366
rect 18256 23344 18552 23364
rect 21256 23420 21552 23440
rect 21312 23418 21336 23420
rect 21392 23418 21416 23420
rect 21472 23418 21496 23420
rect 21334 23366 21336 23418
rect 21398 23366 21410 23418
rect 21472 23366 21474 23418
rect 21312 23364 21336 23366
rect 21392 23364 21416 23366
rect 21472 23364 21496 23366
rect 21256 23344 21552 23364
rect 1756 22876 2052 22896
rect 1812 22874 1836 22876
rect 1892 22874 1916 22876
rect 1972 22874 1996 22876
rect 1834 22822 1836 22874
rect 1898 22822 1910 22874
rect 1972 22822 1974 22874
rect 1812 22820 1836 22822
rect 1892 22820 1916 22822
rect 1972 22820 1996 22822
rect 1756 22800 2052 22820
rect 4756 22876 5052 22896
rect 4812 22874 4836 22876
rect 4892 22874 4916 22876
rect 4972 22874 4996 22876
rect 4834 22822 4836 22874
rect 4898 22822 4910 22874
rect 4972 22822 4974 22874
rect 4812 22820 4836 22822
rect 4892 22820 4916 22822
rect 4972 22820 4996 22822
rect 4756 22800 5052 22820
rect 7756 22876 8052 22896
rect 7812 22874 7836 22876
rect 7892 22874 7916 22876
rect 7972 22874 7996 22876
rect 7834 22822 7836 22874
rect 7898 22822 7910 22874
rect 7972 22822 7974 22874
rect 7812 22820 7836 22822
rect 7892 22820 7916 22822
rect 7972 22820 7996 22822
rect 7756 22800 8052 22820
rect 10756 22876 11052 22896
rect 10812 22874 10836 22876
rect 10892 22874 10916 22876
rect 10972 22874 10996 22876
rect 10834 22822 10836 22874
rect 10898 22822 10910 22874
rect 10972 22822 10974 22874
rect 10812 22820 10836 22822
rect 10892 22820 10916 22822
rect 10972 22820 10996 22822
rect 10756 22800 11052 22820
rect 13756 22876 14052 22896
rect 13812 22874 13836 22876
rect 13892 22874 13916 22876
rect 13972 22874 13996 22876
rect 13834 22822 13836 22874
rect 13898 22822 13910 22874
rect 13972 22822 13974 22874
rect 13812 22820 13836 22822
rect 13892 22820 13916 22822
rect 13972 22820 13996 22822
rect 13756 22800 14052 22820
rect 16756 22876 17052 22896
rect 16812 22874 16836 22876
rect 16892 22874 16916 22876
rect 16972 22874 16996 22876
rect 16834 22822 16836 22874
rect 16898 22822 16910 22874
rect 16972 22822 16974 22874
rect 16812 22820 16836 22822
rect 16892 22820 16916 22822
rect 16972 22820 16996 22822
rect 16756 22800 17052 22820
rect 19756 22876 20052 22896
rect 19812 22874 19836 22876
rect 19892 22874 19916 22876
rect 19972 22874 19996 22876
rect 19834 22822 19836 22874
rect 19898 22822 19910 22874
rect 19972 22822 19974 22874
rect 19812 22820 19836 22822
rect 19892 22820 19916 22822
rect 19972 22820 19996 22822
rect 19756 22800 20052 22820
rect 3256 22332 3552 22352
rect 3312 22330 3336 22332
rect 3392 22330 3416 22332
rect 3472 22330 3496 22332
rect 3334 22278 3336 22330
rect 3398 22278 3410 22330
rect 3472 22278 3474 22330
rect 3312 22276 3336 22278
rect 3392 22276 3416 22278
rect 3472 22276 3496 22278
rect 3256 22256 3552 22276
rect 6256 22332 6552 22352
rect 6312 22330 6336 22332
rect 6392 22330 6416 22332
rect 6472 22330 6496 22332
rect 6334 22278 6336 22330
rect 6398 22278 6410 22330
rect 6472 22278 6474 22330
rect 6312 22276 6336 22278
rect 6392 22276 6416 22278
rect 6472 22276 6496 22278
rect 6256 22256 6552 22276
rect 9256 22332 9552 22352
rect 9312 22330 9336 22332
rect 9392 22330 9416 22332
rect 9472 22330 9496 22332
rect 9334 22278 9336 22330
rect 9398 22278 9410 22330
rect 9472 22278 9474 22330
rect 9312 22276 9336 22278
rect 9392 22276 9416 22278
rect 9472 22276 9496 22278
rect 9256 22256 9552 22276
rect 12256 22332 12552 22352
rect 12312 22330 12336 22332
rect 12392 22330 12416 22332
rect 12472 22330 12496 22332
rect 12334 22278 12336 22330
rect 12398 22278 12410 22330
rect 12472 22278 12474 22330
rect 12312 22276 12336 22278
rect 12392 22276 12416 22278
rect 12472 22276 12496 22278
rect 12256 22256 12552 22276
rect 15256 22332 15552 22352
rect 15312 22330 15336 22332
rect 15392 22330 15416 22332
rect 15472 22330 15496 22332
rect 15334 22278 15336 22330
rect 15398 22278 15410 22330
rect 15472 22278 15474 22330
rect 15312 22276 15336 22278
rect 15392 22276 15416 22278
rect 15472 22276 15496 22278
rect 15256 22256 15552 22276
rect 18256 22332 18552 22352
rect 18312 22330 18336 22332
rect 18392 22330 18416 22332
rect 18472 22330 18496 22332
rect 18334 22278 18336 22330
rect 18398 22278 18410 22330
rect 18472 22278 18474 22330
rect 18312 22276 18336 22278
rect 18392 22276 18416 22278
rect 18472 22276 18496 22278
rect 18256 22256 18552 22276
rect 21256 22332 21552 22352
rect 21312 22330 21336 22332
rect 21392 22330 21416 22332
rect 21472 22330 21496 22332
rect 21334 22278 21336 22330
rect 21398 22278 21410 22330
rect 21472 22278 21474 22330
rect 21312 22276 21336 22278
rect 21392 22276 21416 22278
rect 21472 22276 21496 22278
rect 21256 22256 21552 22276
rect 1756 21788 2052 21808
rect 1812 21786 1836 21788
rect 1892 21786 1916 21788
rect 1972 21786 1996 21788
rect 1834 21734 1836 21786
rect 1898 21734 1910 21786
rect 1972 21734 1974 21786
rect 1812 21732 1836 21734
rect 1892 21732 1916 21734
rect 1972 21732 1996 21734
rect 1756 21712 2052 21732
rect 4756 21788 5052 21808
rect 4812 21786 4836 21788
rect 4892 21786 4916 21788
rect 4972 21786 4996 21788
rect 4834 21734 4836 21786
rect 4898 21734 4910 21786
rect 4972 21734 4974 21786
rect 4812 21732 4836 21734
rect 4892 21732 4916 21734
rect 4972 21732 4996 21734
rect 4756 21712 5052 21732
rect 7756 21788 8052 21808
rect 7812 21786 7836 21788
rect 7892 21786 7916 21788
rect 7972 21786 7996 21788
rect 7834 21734 7836 21786
rect 7898 21734 7910 21786
rect 7972 21734 7974 21786
rect 7812 21732 7836 21734
rect 7892 21732 7916 21734
rect 7972 21732 7996 21734
rect 7756 21712 8052 21732
rect 10756 21788 11052 21808
rect 10812 21786 10836 21788
rect 10892 21786 10916 21788
rect 10972 21786 10996 21788
rect 10834 21734 10836 21786
rect 10898 21734 10910 21786
rect 10972 21734 10974 21786
rect 10812 21732 10836 21734
rect 10892 21732 10916 21734
rect 10972 21732 10996 21734
rect 10756 21712 11052 21732
rect 13756 21788 14052 21808
rect 13812 21786 13836 21788
rect 13892 21786 13916 21788
rect 13972 21786 13996 21788
rect 13834 21734 13836 21786
rect 13898 21734 13910 21786
rect 13972 21734 13974 21786
rect 13812 21732 13836 21734
rect 13892 21732 13916 21734
rect 13972 21732 13996 21734
rect 13756 21712 14052 21732
rect 16756 21788 17052 21808
rect 16812 21786 16836 21788
rect 16892 21786 16916 21788
rect 16972 21786 16996 21788
rect 16834 21734 16836 21786
rect 16898 21734 16910 21786
rect 16972 21734 16974 21786
rect 16812 21732 16836 21734
rect 16892 21732 16916 21734
rect 16972 21732 16996 21734
rect 16756 21712 17052 21732
rect 19756 21788 20052 21808
rect 19812 21786 19836 21788
rect 19892 21786 19916 21788
rect 19972 21786 19996 21788
rect 19834 21734 19836 21786
rect 19898 21734 19910 21786
rect 19972 21734 19974 21786
rect 19812 21732 19836 21734
rect 19892 21732 19916 21734
rect 19972 21732 19996 21734
rect 19756 21712 20052 21732
rect 3256 21244 3552 21264
rect 3312 21242 3336 21244
rect 3392 21242 3416 21244
rect 3472 21242 3496 21244
rect 3334 21190 3336 21242
rect 3398 21190 3410 21242
rect 3472 21190 3474 21242
rect 3312 21188 3336 21190
rect 3392 21188 3416 21190
rect 3472 21188 3496 21190
rect 3256 21168 3552 21188
rect 6256 21244 6552 21264
rect 6312 21242 6336 21244
rect 6392 21242 6416 21244
rect 6472 21242 6496 21244
rect 6334 21190 6336 21242
rect 6398 21190 6410 21242
rect 6472 21190 6474 21242
rect 6312 21188 6336 21190
rect 6392 21188 6416 21190
rect 6472 21188 6496 21190
rect 6256 21168 6552 21188
rect 9256 21244 9552 21264
rect 9312 21242 9336 21244
rect 9392 21242 9416 21244
rect 9472 21242 9496 21244
rect 9334 21190 9336 21242
rect 9398 21190 9410 21242
rect 9472 21190 9474 21242
rect 9312 21188 9336 21190
rect 9392 21188 9416 21190
rect 9472 21188 9496 21190
rect 9256 21168 9552 21188
rect 12256 21244 12552 21264
rect 12312 21242 12336 21244
rect 12392 21242 12416 21244
rect 12472 21242 12496 21244
rect 12334 21190 12336 21242
rect 12398 21190 12410 21242
rect 12472 21190 12474 21242
rect 12312 21188 12336 21190
rect 12392 21188 12416 21190
rect 12472 21188 12496 21190
rect 12256 21168 12552 21188
rect 15256 21244 15552 21264
rect 15312 21242 15336 21244
rect 15392 21242 15416 21244
rect 15472 21242 15496 21244
rect 15334 21190 15336 21242
rect 15398 21190 15410 21242
rect 15472 21190 15474 21242
rect 15312 21188 15336 21190
rect 15392 21188 15416 21190
rect 15472 21188 15496 21190
rect 15256 21168 15552 21188
rect 18256 21244 18552 21264
rect 18312 21242 18336 21244
rect 18392 21242 18416 21244
rect 18472 21242 18496 21244
rect 18334 21190 18336 21242
rect 18398 21190 18410 21242
rect 18472 21190 18474 21242
rect 18312 21188 18336 21190
rect 18392 21188 18416 21190
rect 18472 21188 18496 21190
rect 18256 21168 18552 21188
rect 21256 21244 21552 21264
rect 21312 21242 21336 21244
rect 21392 21242 21416 21244
rect 21472 21242 21496 21244
rect 21334 21190 21336 21242
rect 21398 21190 21410 21242
rect 21472 21190 21474 21242
rect 21312 21188 21336 21190
rect 21392 21188 21416 21190
rect 21472 21188 21496 21190
rect 21256 21168 21552 21188
rect 1756 20700 2052 20720
rect 1812 20698 1836 20700
rect 1892 20698 1916 20700
rect 1972 20698 1996 20700
rect 1834 20646 1836 20698
rect 1898 20646 1910 20698
rect 1972 20646 1974 20698
rect 1812 20644 1836 20646
rect 1892 20644 1916 20646
rect 1972 20644 1996 20646
rect 1756 20624 2052 20644
rect 4756 20700 5052 20720
rect 4812 20698 4836 20700
rect 4892 20698 4916 20700
rect 4972 20698 4996 20700
rect 4834 20646 4836 20698
rect 4898 20646 4910 20698
rect 4972 20646 4974 20698
rect 4812 20644 4836 20646
rect 4892 20644 4916 20646
rect 4972 20644 4996 20646
rect 4756 20624 5052 20644
rect 7756 20700 8052 20720
rect 7812 20698 7836 20700
rect 7892 20698 7916 20700
rect 7972 20698 7996 20700
rect 7834 20646 7836 20698
rect 7898 20646 7910 20698
rect 7972 20646 7974 20698
rect 7812 20644 7836 20646
rect 7892 20644 7916 20646
rect 7972 20644 7996 20646
rect 7756 20624 8052 20644
rect 10756 20700 11052 20720
rect 10812 20698 10836 20700
rect 10892 20698 10916 20700
rect 10972 20698 10996 20700
rect 10834 20646 10836 20698
rect 10898 20646 10910 20698
rect 10972 20646 10974 20698
rect 10812 20644 10836 20646
rect 10892 20644 10916 20646
rect 10972 20644 10996 20646
rect 10756 20624 11052 20644
rect 13756 20700 14052 20720
rect 13812 20698 13836 20700
rect 13892 20698 13916 20700
rect 13972 20698 13996 20700
rect 13834 20646 13836 20698
rect 13898 20646 13910 20698
rect 13972 20646 13974 20698
rect 13812 20644 13836 20646
rect 13892 20644 13916 20646
rect 13972 20644 13996 20646
rect 13756 20624 14052 20644
rect 16756 20700 17052 20720
rect 16812 20698 16836 20700
rect 16892 20698 16916 20700
rect 16972 20698 16996 20700
rect 16834 20646 16836 20698
rect 16898 20646 16910 20698
rect 16972 20646 16974 20698
rect 16812 20644 16836 20646
rect 16892 20644 16916 20646
rect 16972 20644 16996 20646
rect 16756 20624 17052 20644
rect 19756 20700 20052 20720
rect 19812 20698 19836 20700
rect 19892 20698 19916 20700
rect 19972 20698 19996 20700
rect 19834 20646 19836 20698
rect 19898 20646 19910 20698
rect 19972 20646 19974 20698
rect 19812 20644 19836 20646
rect 19892 20644 19916 20646
rect 19972 20644 19996 20646
rect 19756 20624 20052 20644
rect 3256 20156 3552 20176
rect 3312 20154 3336 20156
rect 3392 20154 3416 20156
rect 3472 20154 3496 20156
rect 3334 20102 3336 20154
rect 3398 20102 3410 20154
rect 3472 20102 3474 20154
rect 3312 20100 3336 20102
rect 3392 20100 3416 20102
rect 3472 20100 3496 20102
rect 3256 20080 3552 20100
rect 6256 20156 6552 20176
rect 6312 20154 6336 20156
rect 6392 20154 6416 20156
rect 6472 20154 6496 20156
rect 6334 20102 6336 20154
rect 6398 20102 6410 20154
rect 6472 20102 6474 20154
rect 6312 20100 6336 20102
rect 6392 20100 6416 20102
rect 6472 20100 6496 20102
rect 6256 20080 6552 20100
rect 9256 20156 9552 20176
rect 9312 20154 9336 20156
rect 9392 20154 9416 20156
rect 9472 20154 9496 20156
rect 9334 20102 9336 20154
rect 9398 20102 9410 20154
rect 9472 20102 9474 20154
rect 9312 20100 9336 20102
rect 9392 20100 9416 20102
rect 9472 20100 9496 20102
rect 9256 20080 9552 20100
rect 12256 20156 12552 20176
rect 12312 20154 12336 20156
rect 12392 20154 12416 20156
rect 12472 20154 12496 20156
rect 12334 20102 12336 20154
rect 12398 20102 12410 20154
rect 12472 20102 12474 20154
rect 12312 20100 12336 20102
rect 12392 20100 12416 20102
rect 12472 20100 12496 20102
rect 12256 20080 12552 20100
rect 15256 20156 15552 20176
rect 15312 20154 15336 20156
rect 15392 20154 15416 20156
rect 15472 20154 15496 20156
rect 15334 20102 15336 20154
rect 15398 20102 15410 20154
rect 15472 20102 15474 20154
rect 15312 20100 15336 20102
rect 15392 20100 15416 20102
rect 15472 20100 15496 20102
rect 15256 20080 15552 20100
rect 18256 20156 18552 20176
rect 18312 20154 18336 20156
rect 18392 20154 18416 20156
rect 18472 20154 18496 20156
rect 18334 20102 18336 20154
rect 18398 20102 18410 20154
rect 18472 20102 18474 20154
rect 18312 20100 18336 20102
rect 18392 20100 18416 20102
rect 18472 20100 18496 20102
rect 18256 20080 18552 20100
rect 21256 20156 21552 20176
rect 21312 20154 21336 20156
rect 21392 20154 21416 20156
rect 21472 20154 21496 20156
rect 21334 20102 21336 20154
rect 21398 20102 21410 20154
rect 21472 20102 21474 20154
rect 21312 20100 21336 20102
rect 21392 20100 21416 20102
rect 21472 20100 21496 20102
rect 21256 20080 21552 20100
rect 1756 19612 2052 19632
rect 1812 19610 1836 19612
rect 1892 19610 1916 19612
rect 1972 19610 1996 19612
rect 1834 19558 1836 19610
rect 1898 19558 1910 19610
rect 1972 19558 1974 19610
rect 1812 19556 1836 19558
rect 1892 19556 1916 19558
rect 1972 19556 1996 19558
rect 1756 19536 2052 19556
rect 4756 19612 5052 19632
rect 4812 19610 4836 19612
rect 4892 19610 4916 19612
rect 4972 19610 4996 19612
rect 4834 19558 4836 19610
rect 4898 19558 4910 19610
rect 4972 19558 4974 19610
rect 4812 19556 4836 19558
rect 4892 19556 4916 19558
rect 4972 19556 4996 19558
rect 4756 19536 5052 19556
rect 7756 19612 8052 19632
rect 7812 19610 7836 19612
rect 7892 19610 7916 19612
rect 7972 19610 7996 19612
rect 7834 19558 7836 19610
rect 7898 19558 7910 19610
rect 7972 19558 7974 19610
rect 7812 19556 7836 19558
rect 7892 19556 7916 19558
rect 7972 19556 7996 19558
rect 7756 19536 8052 19556
rect 10756 19612 11052 19632
rect 10812 19610 10836 19612
rect 10892 19610 10916 19612
rect 10972 19610 10996 19612
rect 10834 19558 10836 19610
rect 10898 19558 10910 19610
rect 10972 19558 10974 19610
rect 10812 19556 10836 19558
rect 10892 19556 10916 19558
rect 10972 19556 10996 19558
rect 10756 19536 11052 19556
rect 13756 19612 14052 19632
rect 13812 19610 13836 19612
rect 13892 19610 13916 19612
rect 13972 19610 13996 19612
rect 13834 19558 13836 19610
rect 13898 19558 13910 19610
rect 13972 19558 13974 19610
rect 13812 19556 13836 19558
rect 13892 19556 13916 19558
rect 13972 19556 13996 19558
rect 13756 19536 14052 19556
rect 16756 19612 17052 19632
rect 16812 19610 16836 19612
rect 16892 19610 16916 19612
rect 16972 19610 16996 19612
rect 16834 19558 16836 19610
rect 16898 19558 16910 19610
rect 16972 19558 16974 19610
rect 16812 19556 16836 19558
rect 16892 19556 16916 19558
rect 16972 19556 16996 19558
rect 16756 19536 17052 19556
rect 19756 19612 20052 19632
rect 19812 19610 19836 19612
rect 19892 19610 19916 19612
rect 19972 19610 19996 19612
rect 19834 19558 19836 19610
rect 19898 19558 19910 19610
rect 19972 19558 19974 19610
rect 19812 19556 19836 19558
rect 19892 19556 19916 19558
rect 19972 19556 19996 19558
rect 19756 19536 20052 19556
rect 3256 19068 3552 19088
rect 3312 19066 3336 19068
rect 3392 19066 3416 19068
rect 3472 19066 3496 19068
rect 3334 19014 3336 19066
rect 3398 19014 3410 19066
rect 3472 19014 3474 19066
rect 3312 19012 3336 19014
rect 3392 19012 3416 19014
rect 3472 19012 3496 19014
rect 3256 18992 3552 19012
rect 6256 19068 6552 19088
rect 6312 19066 6336 19068
rect 6392 19066 6416 19068
rect 6472 19066 6496 19068
rect 6334 19014 6336 19066
rect 6398 19014 6410 19066
rect 6472 19014 6474 19066
rect 6312 19012 6336 19014
rect 6392 19012 6416 19014
rect 6472 19012 6496 19014
rect 6256 18992 6552 19012
rect 9256 19068 9552 19088
rect 9312 19066 9336 19068
rect 9392 19066 9416 19068
rect 9472 19066 9496 19068
rect 9334 19014 9336 19066
rect 9398 19014 9410 19066
rect 9472 19014 9474 19066
rect 9312 19012 9336 19014
rect 9392 19012 9416 19014
rect 9472 19012 9496 19014
rect 9256 18992 9552 19012
rect 12256 19068 12552 19088
rect 12312 19066 12336 19068
rect 12392 19066 12416 19068
rect 12472 19066 12496 19068
rect 12334 19014 12336 19066
rect 12398 19014 12410 19066
rect 12472 19014 12474 19066
rect 12312 19012 12336 19014
rect 12392 19012 12416 19014
rect 12472 19012 12496 19014
rect 12256 18992 12552 19012
rect 15256 19068 15552 19088
rect 15312 19066 15336 19068
rect 15392 19066 15416 19068
rect 15472 19066 15496 19068
rect 15334 19014 15336 19066
rect 15398 19014 15410 19066
rect 15472 19014 15474 19066
rect 15312 19012 15336 19014
rect 15392 19012 15416 19014
rect 15472 19012 15496 19014
rect 15256 18992 15552 19012
rect 18256 19068 18552 19088
rect 18312 19066 18336 19068
rect 18392 19066 18416 19068
rect 18472 19066 18496 19068
rect 18334 19014 18336 19066
rect 18398 19014 18410 19066
rect 18472 19014 18474 19066
rect 18312 19012 18336 19014
rect 18392 19012 18416 19014
rect 18472 19012 18496 19014
rect 18256 18992 18552 19012
rect 21256 19068 21552 19088
rect 21312 19066 21336 19068
rect 21392 19066 21416 19068
rect 21472 19066 21496 19068
rect 21334 19014 21336 19066
rect 21398 19014 21410 19066
rect 21472 19014 21474 19066
rect 21312 19012 21336 19014
rect 21392 19012 21416 19014
rect 21472 19012 21496 19014
rect 21256 18992 21552 19012
rect 1756 18524 2052 18544
rect 1812 18522 1836 18524
rect 1892 18522 1916 18524
rect 1972 18522 1996 18524
rect 1834 18470 1836 18522
rect 1898 18470 1910 18522
rect 1972 18470 1974 18522
rect 1812 18468 1836 18470
rect 1892 18468 1916 18470
rect 1972 18468 1996 18470
rect 1756 18448 2052 18468
rect 4756 18524 5052 18544
rect 4812 18522 4836 18524
rect 4892 18522 4916 18524
rect 4972 18522 4996 18524
rect 4834 18470 4836 18522
rect 4898 18470 4910 18522
rect 4972 18470 4974 18522
rect 4812 18468 4836 18470
rect 4892 18468 4916 18470
rect 4972 18468 4996 18470
rect 4756 18448 5052 18468
rect 7756 18524 8052 18544
rect 7812 18522 7836 18524
rect 7892 18522 7916 18524
rect 7972 18522 7996 18524
rect 7834 18470 7836 18522
rect 7898 18470 7910 18522
rect 7972 18470 7974 18522
rect 7812 18468 7836 18470
rect 7892 18468 7916 18470
rect 7972 18468 7996 18470
rect 7756 18448 8052 18468
rect 10756 18524 11052 18544
rect 10812 18522 10836 18524
rect 10892 18522 10916 18524
rect 10972 18522 10996 18524
rect 10834 18470 10836 18522
rect 10898 18470 10910 18522
rect 10972 18470 10974 18522
rect 10812 18468 10836 18470
rect 10892 18468 10916 18470
rect 10972 18468 10996 18470
rect 10756 18448 11052 18468
rect 13756 18524 14052 18544
rect 13812 18522 13836 18524
rect 13892 18522 13916 18524
rect 13972 18522 13996 18524
rect 13834 18470 13836 18522
rect 13898 18470 13910 18522
rect 13972 18470 13974 18522
rect 13812 18468 13836 18470
rect 13892 18468 13916 18470
rect 13972 18468 13996 18470
rect 13756 18448 14052 18468
rect 16756 18524 17052 18544
rect 16812 18522 16836 18524
rect 16892 18522 16916 18524
rect 16972 18522 16996 18524
rect 16834 18470 16836 18522
rect 16898 18470 16910 18522
rect 16972 18470 16974 18522
rect 16812 18468 16836 18470
rect 16892 18468 16916 18470
rect 16972 18468 16996 18470
rect 16756 18448 17052 18468
rect 19756 18524 20052 18544
rect 19812 18522 19836 18524
rect 19892 18522 19916 18524
rect 19972 18522 19996 18524
rect 19834 18470 19836 18522
rect 19898 18470 19910 18522
rect 19972 18470 19974 18522
rect 19812 18468 19836 18470
rect 19892 18468 19916 18470
rect 19972 18468 19996 18470
rect 19756 18448 20052 18468
rect 3256 17980 3552 18000
rect 3312 17978 3336 17980
rect 3392 17978 3416 17980
rect 3472 17978 3496 17980
rect 3334 17926 3336 17978
rect 3398 17926 3410 17978
rect 3472 17926 3474 17978
rect 3312 17924 3336 17926
rect 3392 17924 3416 17926
rect 3472 17924 3496 17926
rect 3256 17904 3552 17924
rect 6256 17980 6552 18000
rect 6312 17978 6336 17980
rect 6392 17978 6416 17980
rect 6472 17978 6496 17980
rect 6334 17926 6336 17978
rect 6398 17926 6410 17978
rect 6472 17926 6474 17978
rect 6312 17924 6336 17926
rect 6392 17924 6416 17926
rect 6472 17924 6496 17926
rect 6256 17904 6552 17924
rect 9256 17980 9552 18000
rect 9312 17978 9336 17980
rect 9392 17978 9416 17980
rect 9472 17978 9496 17980
rect 9334 17926 9336 17978
rect 9398 17926 9410 17978
rect 9472 17926 9474 17978
rect 9312 17924 9336 17926
rect 9392 17924 9416 17926
rect 9472 17924 9496 17926
rect 9256 17904 9552 17924
rect 12256 17980 12552 18000
rect 12312 17978 12336 17980
rect 12392 17978 12416 17980
rect 12472 17978 12496 17980
rect 12334 17926 12336 17978
rect 12398 17926 12410 17978
rect 12472 17926 12474 17978
rect 12312 17924 12336 17926
rect 12392 17924 12416 17926
rect 12472 17924 12496 17926
rect 12256 17904 12552 17924
rect 15256 17980 15552 18000
rect 15312 17978 15336 17980
rect 15392 17978 15416 17980
rect 15472 17978 15496 17980
rect 15334 17926 15336 17978
rect 15398 17926 15410 17978
rect 15472 17926 15474 17978
rect 15312 17924 15336 17926
rect 15392 17924 15416 17926
rect 15472 17924 15496 17926
rect 15256 17904 15552 17924
rect 18256 17980 18552 18000
rect 18312 17978 18336 17980
rect 18392 17978 18416 17980
rect 18472 17978 18496 17980
rect 18334 17926 18336 17978
rect 18398 17926 18410 17978
rect 18472 17926 18474 17978
rect 18312 17924 18336 17926
rect 18392 17924 18416 17926
rect 18472 17924 18496 17926
rect 18256 17904 18552 17924
rect 21256 17980 21552 18000
rect 21312 17978 21336 17980
rect 21392 17978 21416 17980
rect 21472 17978 21496 17980
rect 21334 17926 21336 17978
rect 21398 17926 21410 17978
rect 21472 17926 21474 17978
rect 21312 17924 21336 17926
rect 21392 17924 21416 17926
rect 21472 17924 21496 17926
rect 21256 17904 21552 17924
rect 1756 17436 2052 17456
rect 1812 17434 1836 17436
rect 1892 17434 1916 17436
rect 1972 17434 1996 17436
rect 1834 17382 1836 17434
rect 1898 17382 1910 17434
rect 1972 17382 1974 17434
rect 1812 17380 1836 17382
rect 1892 17380 1916 17382
rect 1972 17380 1996 17382
rect 1756 17360 2052 17380
rect 4756 17436 5052 17456
rect 4812 17434 4836 17436
rect 4892 17434 4916 17436
rect 4972 17434 4996 17436
rect 4834 17382 4836 17434
rect 4898 17382 4910 17434
rect 4972 17382 4974 17434
rect 4812 17380 4836 17382
rect 4892 17380 4916 17382
rect 4972 17380 4996 17382
rect 4756 17360 5052 17380
rect 7756 17436 8052 17456
rect 7812 17434 7836 17436
rect 7892 17434 7916 17436
rect 7972 17434 7996 17436
rect 7834 17382 7836 17434
rect 7898 17382 7910 17434
rect 7972 17382 7974 17434
rect 7812 17380 7836 17382
rect 7892 17380 7916 17382
rect 7972 17380 7996 17382
rect 7756 17360 8052 17380
rect 10756 17436 11052 17456
rect 10812 17434 10836 17436
rect 10892 17434 10916 17436
rect 10972 17434 10996 17436
rect 10834 17382 10836 17434
rect 10898 17382 10910 17434
rect 10972 17382 10974 17434
rect 10812 17380 10836 17382
rect 10892 17380 10916 17382
rect 10972 17380 10996 17382
rect 10756 17360 11052 17380
rect 13756 17436 14052 17456
rect 13812 17434 13836 17436
rect 13892 17434 13916 17436
rect 13972 17434 13996 17436
rect 13834 17382 13836 17434
rect 13898 17382 13910 17434
rect 13972 17382 13974 17434
rect 13812 17380 13836 17382
rect 13892 17380 13916 17382
rect 13972 17380 13996 17382
rect 13756 17360 14052 17380
rect 16756 17436 17052 17456
rect 16812 17434 16836 17436
rect 16892 17434 16916 17436
rect 16972 17434 16996 17436
rect 16834 17382 16836 17434
rect 16898 17382 16910 17434
rect 16972 17382 16974 17434
rect 16812 17380 16836 17382
rect 16892 17380 16916 17382
rect 16972 17380 16996 17382
rect 16756 17360 17052 17380
rect 19756 17436 20052 17456
rect 19812 17434 19836 17436
rect 19892 17434 19916 17436
rect 19972 17434 19996 17436
rect 19834 17382 19836 17434
rect 19898 17382 19910 17434
rect 19972 17382 19974 17434
rect 19812 17380 19836 17382
rect 19892 17380 19916 17382
rect 19972 17380 19996 17382
rect 19756 17360 20052 17380
rect 3256 16892 3552 16912
rect 3312 16890 3336 16892
rect 3392 16890 3416 16892
rect 3472 16890 3496 16892
rect 3334 16838 3336 16890
rect 3398 16838 3410 16890
rect 3472 16838 3474 16890
rect 3312 16836 3336 16838
rect 3392 16836 3416 16838
rect 3472 16836 3496 16838
rect 3256 16816 3552 16836
rect 6256 16892 6552 16912
rect 6312 16890 6336 16892
rect 6392 16890 6416 16892
rect 6472 16890 6496 16892
rect 6334 16838 6336 16890
rect 6398 16838 6410 16890
rect 6472 16838 6474 16890
rect 6312 16836 6336 16838
rect 6392 16836 6416 16838
rect 6472 16836 6496 16838
rect 6256 16816 6552 16836
rect 9256 16892 9552 16912
rect 9312 16890 9336 16892
rect 9392 16890 9416 16892
rect 9472 16890 9496 16892
rect 9334 16838 9336 16890
rect 9398 16838 9410 16890
rect 9472 16838 9474 16890
rect 9312 16836 9336 16838
rect 9392 16836 9416 16838
rect 9472 16836 9496 16838
rect 9256 16816 9552 16836
rect 12256 16892 12552 16912
rect 12312 16890 12336 16892
rect 12392 16890 12416 16892
rect 12472 16890 12496 16892
rect 12334 16838 12336 16890
rect 12398 16838 12410 16890
rect 12472 16838 12474 16890
rect 12312 16836 12336 16838
rect 12392 16836 12416 16838
rect 12472 16836 12496 16838
rect 12256 16816 12552 16836
rect 15256 16892 15552 16912
rect 15312 16890 15336 16892
rect 15392 16890 15416 16892
rect 15472 16890 15496 16892
rect 15334 16838 15336 16890
rect 15398 16838 15410 16890
rect 15472 16838 15474 16890
rect 15312 16836 15336 16838
rect 15392 16836 15416 16838
rect 15472 16836 15496 16838
rect 15256 16816 15552 16836
rect 18256 16892 18552 16912
rect 18312 16890 18336 16892
rect 18392 16890 18416 16892
rect 18472 16890 18496 16892
rect 18334 16838 18336 16890
rect 18398 16838 18410 16890
rect 18472 16838 18474 16890
rect 18312 16836 18336 16838
rect 18392 16836 18416 16838
rect 18472 16836 18496 16838
rect 18256 16816 18552 16836
rect 21256 16892 21552 16912
rect 21312 16890 21336 16892
rect 21392 16890 21416 16892
rect 21472 16890 21496 16892
rect 21334 16838 21336 16890
rect 21398 16838 21410 16890
rect 21472 16838 21474 16890
rect 21312 16836 21336 16838
rect 21392 16836 21416 16838
rect 21472 16836 21496 16838
rect 21256 16816 21552 16836
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 1756 16348 2052 16368
rect 1812 16346 1836 16348
rect 1892 16346 1916 16348
rect 1972 16346 1996 16348
rect 1834 16294 1836 16346
rect 1898 16294 1910 16346
rect 1972 16294 1974 16346
rect 1812 16292 1836 16294
rect 1892 16292 1916 16294
rect 1972 16292 1996 16294
rect 1756 16272 2052 16292
rect 4756 16348 5052 16368
rect 4812 16346 4836 16348
rect 4892 16346 4916 16348
rect 4972 16346 4996 16348
rect 4834 16294 4836 16346
rect 4898 16294 4910 16346
rect 4972 16294 4974 16346
rect 4812 16292 4836 16294
rect 4892 16292 4916 16294
rect 4972 16292 4996 16294
rect 4756 16272 5052 16292
rect 7756 16348 8052 16368
rect 7812 16346 7836 16348
rect 7892 16346 7916 16348
rect 7972 16346 7996 16348
rect 7834 16294 7836 16346
rect 7898 16294 7910 16346
rect 7972 16294 7974 16346
rect 7812 16292 7836 16294
rect 7892 16292 7916 16294
rect 7972 16292 7996 16294
rect 7756 16272 8052 16292
rect 10756 16348 11052 16368
rect 10812 16346 10836 16348
rect 10892 16346 10916 16348
rect 10972 16346 10996 16348
rect 10834 16294 10836 16346
rect 10898 16294 10910 16346
rect 10972 16294 10974 16346
rect 10812 16292 10836 16294
rect 10892 16292 10916 16294
rect 10972 16292 10996 16294
rect 10756 16272 11052 16292
rect 13756 16348 14052 16368
rect 13812 16346 13836 16348
rect 13892 16346 13916 16348
rect 13972 16346 13996 16348
rect 13834 16294 13836 16346
rect 13898 16294 13910 16346
rect 13972 16294 13974 16346
rect 13812 16292 13836 16294
rect 13892 16292 13916 16294
rect 13972 16292 13996 16294
rect 13756 16272 14052 16292
rect 14108 15910 14136 16526
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 3256 15804 3552 15824
rect 3312 15802 3336 15804
rect 3392 15802 3416 15804
rect 3472 15802 3496 15804
rect 3334 15750 3336 15802
rect 3398 15750 3410 15802
rect 3472 15750 3474 15802
rect 3312 15748 3336 15750
rect 3392 15748 3416 15750
rect 3472 15748 3496 15750
rect 3256 15728 3552 15748
rect 6256 15804 6552 15824
rect 6312 15802 6336 15804
rect 6392 15802 6416 15804
rect 6472 15802 6496 15804
rect 6334 15750 6336 15802
rect 6398 15750 6410 15802
rect 6472 15750 6474 15802
rect 6312 15748 6336 15750
rect 6392 15748 6416 15750
rect 6472 15748 6496 15750
rect 6256 15728 6552 15748
rect 9256 15804 9552 15824
rect 9312 15802 9336 15804
rect 9392 15802 9416 15804
rect 9472 15802 9496 15804
rect 9334 15750 9336 15802
rect 9398 15750 9410 15802
rect 9472 15750 9474 15802
rect 9312 15748 9336 15750
rect 9392 15748 9416 15750
rect 9472 15748 9496 15750
rect 9256 15728 9552 15748
rect 12256 15804 12552 15824
rect 12312 15802 12336 15804
rect 12392 15802 12416 15804
rect 12472 15802 12496 15804
rect 12334 15750 12336 15802
rect 12398 15750 12410 15802
rect 12472 15750 12474 15802
rect 12312 15748 12336 15750
rect 12392 15748 12416 15750
rect 12472 15748 12496 15750
rect 12256 15728 12552 15748
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 1756 15260 2052 15280
rect 1812 15258 1836 15260
rect 1892 15258 1916 15260
rect 1972 15258 1996 15260
rect 1834 15206 1836 15258
rect 1898 15206 1910 15258
rect 1972 15206 1974 15258
rect 1812 15204 1836 15206
rect 1892 15204 1916 15206
rect 1972 15204 1996 15206
rect 1756 15184 2052 15204
rect 4756 15260 5052 15280
rect 4812 15258 4836 15260
rect 4892 15258 4916 15260
rect 4972 15258 4996 15260
rect 4834 15206 4836 15258
rect 4898 15206 4910 15258
rect 4972 15206 4974 15258
rect 4812 15204 4836 15206
rect 4892 15204 4916 15206
rect 4972 15204 4996 15206
rect 4756 15184 5052 15204
rect 7756 15260 8052 15280
rect 7812 15258 7836 15260
rect 7892 15258 7916 15260
rect 7972 15258 7996 15260
rect 7834 15206 7836 15258
rect 7898 15206 7910 15258
rect 7972 15206 7974 15258
rect 7812 15204 7836 15206
rect 7892 15204 7916 15206
rect 7972 15204 7996 15206
rect 7756 15184 8052 15204
rect 10756 15260 11052 15280
rect 10812 15258 10836 15260
rect 10892 15258 10916 15260
rect 10972 15258 10996 15260
rect 10834 15206 10836 15258
rect 10898 15206 10910 15258
rect 10972 15206 10974 15258
rect 10812 15204 10836 15206
rect 10892 15204 10916 15206
rect 10972 15204 10996 15206
rect 10756 15184 11052 15204
rect 12728 15162 12756 15438
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 3256 14716 3552 14736
rect 3312 14714 3336 14716
rect 3392 14714 3416 14716
rect 3472 14714 3496 14716
rect 3334 14662 3336 14714
rect 3398 14662 3410 14714
rect 3472 14662 3474 14714
rect 3312 14660 3336 14662
rect 3392 14660 3416 14662
rect 3472 14660 3496 14662
rect 3256 14640 3552 14660
rect 6256 14716 6552 14736
rect 6312 14714 6336 14716
rect 6392 14714 6416 14716
rect 6472 14714 6496 14716
rect 6334 14662 6336 14714
rect 6398 14662 6410 14714
rect 6472 14662 6474 14714
rect 6312 14660 6336 14662
rect 6392 14660 6416 14662
rect 6472 14660 6496 14662
rect 6256 14640 6552 14660
rect 9256 14716 9552 14736
rect 9312 14714 9336 14716
rect 9392 14714 9416 14716
rect 9472 14714 9496 14716
rect 9334 14662 9336 14714
rect 9398 14662 9410 14714
rect 9472 14662 9474 14714
rect 9312 14660 9336 14662
rect 9392 14660 9416 14662
rect 9472 14660 9496 14662
rect 9256 14640 9552 14660
rect 12256 14716 12552 14736
rect 12312 14714 12336 14716
rect 12392 14714 12416 14716
rect 12472 14714 12496 14716
rect 12334 14662 12336 14714
rect 12398 14662 12410 14714
rect 12472 14662 12474 14714
rect 12312 14660 12336 14662
rect 12392 14660 12416 14662
rect 12472 14660 12496 14662
rect 12256 14640 12552 14660
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 1756 14172 2052 14192
rect 1812 14170 1836 14172
rect 1892 14170 1916 14172
rect 1972 14170 1996 14172
rect 1834 14118 1836 14170
rect 1898 14118 1910 14170
rect 1972 14118 1974 14170
rect 1812 14116 1836 14118
rect 1892 14116 1916 14118
rect 1972 14116 1996 14118
rect 1756 14096 2052 14116
rect 4756 14172 5052 14192
rect 4812 14170 4836 14172
rect 4892 14170 4916 14172
rect 4972 14170 4996 14172
rect 4834 14118 4836 14170
rect 4898 14118 4910 14170
rect 4972 14118 4974 14170
rect 4812 14116 4836 14118
rect 4892 14116 4916 14118
rect 4972 14116 4996 14118
rect 4756 14096 5052 14116
rect 7756 14172 8052 14192
rect 7812 14170 7836 14172
rect 7892 14170 7916 14172
rect 7972 14170 7996 14172
rect 7834 14118 7836 14170
rect 7898 14118 7910 14170
rect 7972 14118 7974 14170
rect 7812 14116 7836 14118
rect 7892 14116 7916 14118
rect 7972 14116 7996 14118
rect 7756 14096 8052 14116
rect 10756 14172 11052 14192
rect 10812 14170 10836 14172
rect 10892 14170 10916 14172
rect 10972 14170 10996 14172
rect 10834 14118 10836 14170
rect 10898 14118 10910 14170
rect 10972 14118 10974 14170
rect 10812 14116 10836 14118
rect 10892 14116 10916 14118
rect 10972 14116 10996 14118
rect 10756 14096 11052 14116
rect 11900 14006 11928 14418
rect 12912 14346 12940 15302
rect 13280 15026 13308 15302
rect 13756 15260 14052 15280
rect 13812 15258 13836 15260
rect 13892 15258 13916 15260
rect 13972 15258 13996 15260
rect 13834 15206 13836 15258
rect 13898 15206 13910 15258
rect 13972 15206 13974 15258
rect 13812 15204 13836 15206
rect 13892 15204 13916 15206
rect 13972 15204 13996 15206
rect 13756 15184 14052 15204
rect 14108 15162 14136 15846
rect 14200 15366 14228 15982
rect 14292 15706 14320 16390
rect 14936 16182 14964 16390
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14556 16040 14608 16046
rect 14608 16000 14688 16028
rect 14556 15982 14608 15988
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14660 15366 14688 16000
rect 15580 15978 15608 16526
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15256 15804 15552 15824
rect 15312 15802 15336 15804
rect 15392 15802 15416 15804
rect 15472 15802 15496 15804
rect 15334 15750 15336 15802
rect 15398 15750 15410 15802
rect 15472 15750 15474 15802
rect 15312 15748 15336 15750
rect 15392 15748 15416 15750
rect 15472 15748 15496 15750
rect 15256 15728 15552 15748
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12176 14074 12204 14282
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 110 13696 166 13705
rect 110 13631 166 13640
rect 124 12209 152 13631
rect 3256 13628 3552 13648
rect 3312 13626 3336 13628
rect 3392 13626 3416 13628
rect 3472 13626 3496 13628
rect 3334 13574 3336 13626
rect 3398 13574 3410 13626
rect 3472 13574 3474 13626
rect 3312 13572 3336 13574
rect 3392 13572 3416 13574
rect 3472 13572 3496 13574
rect 3256 13552 3552 13572
rect 6256 13628 6552 13648
rect 6312 13626 6336 13628
rect 6392 13626 6416 13628
rect 6472 13626 6496 13628
rect 6334 13574 6336 13626
rect 6398 13574 6410 13626
rect 6472 13574 6474 13626
rect 6312 13572 6336 13574
rect 6392 13572 6416 13574
rect 6472 13572 6496 13574
rect 6256 13552 6552 13572
rect 8680 13190 8708 13874
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 9256 13628 9552 13648
rect 9312 13626 9336 13628
rect 9392 13626 9416 13628
rect 9472 13626 9496 13628
rect 9334 13574 9336 13626
rect 9398 13574 9410 13626
rect 9472 13574 9474 13626
rect 9312 13572 9336 13574
rect 9392 13572 9416 13574
rect 9472 13572 9496 13574
rect 9256 13552 9552 13572
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 1756 13084 2052 13104
rect 1812 13082 1836 13084
rect 1892 13082 1916 13084
rect 1972 13082 1996 13084
rect 1834 13030 1836 13082
rect 1898 13030 1910 13082
rect 1972 13030 1974 13082
rect 1812 13028 1836 13030
rect 1892 13028 1916 13030
rect 1972 13028 1996 13030
rect 1756 13008 2052 13028
rect 4756 13084 5052 13104
rect 4812 13082 4836 13084
rect 4892 13082 4916 13084
rect 4972 13082 4996 13084
rect 4834 13030 4836 13082
rect 4898 13030 4910 13082
rect 4972 13030 4974 13082
rect 4812 13028 4836 13030
rect 4892 13028 4916 13030
rect 4972 13028 4996 13030
rect 4756 13008 5052 13028
rect 7756 13084 8052 13104
rect 7812 13082 7836 13084
rect 7892 13082 7916 13084
rect 7972 13082 7996 13084
rect 7834 13030 7836 13082
rect 7898 13030 7910 13082
rect 7972 13030 7974 13082
rect 7812 13028 7836 13030
rect 7892 13028 7916 13030
rect 7972 13028 7996 13030
rect 7756 13008 8052 13028
rect 3256 12540 3552 12560
rect 3312 12538 3336 12540
rect 3392 12538 3416 12540
rect 3472 12538 3496 12540
rect 3334 12486 3336 12538
rect 3398 12486 3410 12538
rect 3472 12486 3474 12538
rect 3312 12484 3336 12486
rect 3392 12484 3416 12486
rect 3472 12484 3496 12486
rect 3256 12464 3552 12484
rect 6256 12540 6552 12560
rect 6312 12538 6336 12540
rect 6392 12538 6416 12540
rect 6472 12538 6496 12540
rect 6334 12486 6336 12538
rect 6398 12486 6410 12538
rect 6472 12486 6474 12538
rect 6312 12484 6336 12486
rect 6392 12484 6416 12486
rect 6472 12484 6496 12486
rect 6256 12464 6552 12484
rect 8404 12442 8432 13126
rect 10756 13084 11052 13104
rect 10812 13082 10836 13084
rect 10892 13082 10916 13084
rect 10972 13082 10996 13084
rect 10834 13030 10836 13082
rect 10898 13030 10910 13082
rect 10972 13030 10974 13082
rect 10812 13028 10836 13030
rect 10892 13028 10916 13030
rect 10972 13028 10996 13030
rect 10756 13008 11052 13028
rect 11256 12986 11284 13670
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 9256 12540 9552 12560
rect 9312 12538 9336 12540
rect 9392 12538 9416 12540
rect 9472 12538 9496 12540
rect 9334 12486 9336 12538
rect 9398 12486 9410 12538
rect 9472 12486 9474 12538
rect 9312 12484 9336 12486
rect 9392 12484 9416 12486
rect 9472 12484 9496 12486
rect 9256 12464 9552 12484
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 110 12200 166 12209
rect 110 12135 166 12144
rect 1756 11996 2052 12016
rect 1812 11994 1836 11996
rect 1892 11994 1916 11996
rect 1972 11994 1996 11996
rect 1834 11942 1836 11994
rect 1898 11942 1910 11994
rect 1972 11942 1974 11994
rect 1812 11940 1836 11942
rect 1892 11940 1916 11942
rect 1972 11940 1996 11942
rect 1756 11920 2052 11940
rect 4756 11996 5052 12016
rect 4812 11994 4836 11996
rect 4892 11994 4916 11996
rect 4972 11994 4996 11996
rect 4834 11942 4836 11994
rect 4898 11942 4910 11994
rect 4972 11942 4974 11994
rect 4812 11940 4836 11942
rect 4892 11940 4916 11942
rect 4972 11940 4996 11942
rect 4756 11920 5052 11940
rect 7756 11996 8052 12016
rect 7812 11994 7836 11996
rect 7892 11994 7916 11996
rect 7972 11994 7996 11996
rect 7834 11942 7836 11994
rect 7898 11942 7910 11994
rect 7972 11942 7974 11994
rect 7812 11940 7836 11942
rect 7892 11940 7916 11942
rect 7972 11940 7996 11942
rect 7756 11920 8052 11940
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 3256 11452 3552 11472
rect 3312 11450 3336 11452
rect 3392 11450 3416 11452
rect 3472 11450 3496 11452
rect 3334 11398 3336 11450
rect 3398 11398 3410 11450
rect 3472 11398 3474 11450
rect 3312 11396 3336 11398
rect 3392 11396 3416 11398
rect 3472 11396 3496 11398
rect 3256 11376 3552 11396
rect 1756 10908 2052 10928
rect 1812 10906 1836 10908
rect 1892 10906 1916 10908
rect 1972 10906 1996 10908
rect 1834 10854 1836 10906
rect 1898 10854 1910 10906
rect 1972 10854 1974 10906
rect 1812 10852 1836 10854
rect 1892 10852 1916 10854
rect 1972 10852 1996 10854
rect 1756 10832 2052 10852
rect 4756 10908 5052 10928
rect 4812 10906 4836 10908
rect 4892 10906 4916 10908
rect 4972 10906 4996 10908
rect 4834 10854 4836 10906
rect 4898 10854 4910 10906
rect 4972 10854 4974 10906
rect 4812 10852 4836 10854
rect 4892 10852 4916 10854
rect 4972 10852 4996 10854
rect 4756 10832 5052 10852
rect 3256 10364 3552 10384
rect 3312 10362 3336 10364
rect 3392 10362 3416 10364
rect 3472 10362 3496 10364
rect 3334 10310 3336 10362
rect 3398 10310 3410 10362
rect 3472 10310 3474 10362
rect 3312 10308 3336 10310
rect 3392 10308 3416 10310
rect 3472 10308 3496 10310
rect 3256 10288 3552 10308
rect 6196 10062 6224 11494
rect 6256 11452 6552 11472
rect 6312 11450 6336 11452
rect 6392 11450 6416 11452
rect 6472 11450 6496 11452
rect 6334 11398 6336 11450
rect 6398 11398 6410 11450
rect 6472 11398 6474 11450
rect 6312 11396 6336 11398
rect 6392 11396 6416 11398
rect 6472 11396 6496 11398
rect 6256 11376 6552 11396
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10470 6776 11086
rect 8036 11082 8064 11630
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6256 10364 6552 10384
rect 6312 10362 6336 10364
rect 6392 10362 6416 10364
rect 6472 10362 6496 10364
rect 6334 10310 6336 10362
rect 6398 10310 6410 10362
rect 6472 10310 6474 10362
rect 6312 10308 6336 10310
rect 6392 10308 6416 10310
rect 6472 10308 6496 10310
rect 6256 10288 6552 10308
rect 6748 10266 6776 10406
rect 6932 10266 6960 10950
rect 7756 10908 8052 10928
rect 7812 10906 7836 10908
rect 7892 10906 7916 10908
rect 7972 10906 7996 10908
rect 7834 10854 7836 10906
rect 7898 10854 7910 10906
rect 7972 10854 7974 10906
rect 7812 10852 7836 10854
rect 7892 10852 7916 10854
rect 7972 10852 7996 10854
rect 7756 10832 8052 10852
rect 8128 10810 8156 11086
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6932 10062 6960 10202
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 1756 9820 2052 9840
rect 1812 9818 1836 9820
rect 1892 9818 1916 9820
rect 1972 9818 1996 9820
rect 1834 9766 1836 9818
rect 1898 9766 1910 9818
rect 1972 9766 1974 9818
rect 1812 9764 1836 9766
rect 1892 9764 1916 9766
rect 1972 9764 1996 9766
rect 1756 9744 2052 9764
rect 4756 9820 5052 9840
rect 4812 9818 4836 9820
rect 4892 9818 4916 9820
rect 4972 9818 4996 9820
rect 4834 9766 4836 9818
rect 4898 9766 4910 9818
rect 4972 9766 4974 9818
rect 4812 9764 4836 9766
rect 4892 9764 4916 9766
rect 4972 9764 4996 9766
rect 4756 9744 5052 9764
rect 6196 9654 6224 9998
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 7300 9518 7328 9930
rect 7576 9654 7604 9930
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7012 9512 7064 9518
rect 7288 9512 7340 9518
rect 7064 9472 7144 9500
rect 7012 9454 7064 9460
rect 3256 9276 3552 9296
rect 3312 9274 3336 9276
rect 3392 9274 3416 9276
rect 3472 9274 3496 9276
rect 3334 9222 3336 9274
rect 3398 9222 3410 9274
rect 3472 9222 3474 9274
rect 3312 9220 3336 9222
rect 3392 9220 3416 9222
rect 3472 9220 3496 9222
rect 3256 9200 3552 9220
rect 6256 9276 6552 9296
rect 6312 9274 6336 9276
rect 6392 9274 6416 9276
rect 6472 9274 6496 9276
rect 6334 9222 6336 9274
rect 6398 9222 6410 9274
rect 6472 9222 6474 9274
rect 6312 9220 6336 9222
rect 6392 9220 6416 9222
rect 6472 9220 6496 9222
rect 6256 9200 6552 9220
rect 7116 9042 7144 9472
rect 7288 9454 7340 9460
rect 7300 9178 7328 9454
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 1756 8732 2052 8752
rect 1812 8730 1836 8732
rect 1892 8730 1916 8732
rect 1972 8730 1996 8732
rect 1834 8678 1836 8730
rect 1898 8678 1910 8730
rect 1972 8678 1974 8730
rect 1812 8676 1836 8678
rect 1892 8676 1916 8678
rect 1972 8676 1996 8678
rect 1756 8656 2052 8676
rect 4756 8732 5052 8752
rect 4812 8730 4836 8732
rect 4892 8730 4916 8732
rect 4972 8730 4996 8732
rect 4834 8678 4836 8730
rect 4898 8678 4910 8730
rect 4972 8678 4974 8730
rect 4812 8676 4836 8678
rect 4892 8676 4916 8678
rect 4972 8676 4996 8678
rect 4756 8656 5052 8676
rect 6104 8294 6132 8910
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 3256 8188 3552 8208
rect 3312 8186 3336 8188
rect 3392 8186 3416 8188
rect 3472 8186 3496 8188
rect 3334 8134 3336 8186
rect 3398 8134 3410 8186
rect 3472 8134 3474 8186
rect 3312 8132 3336 8134
rect 3392 8132 3416 8134
rect 3472 8132 3496 8134
rect 3256 8112 3552 8132
rect 1756 7644 2052 7664
rect 1812 7642 1836 7644
rect 1892 7642 1916 7644
rect 1972 7642 1996 7644
rect 1834 7590 1836 7642
rect 1898 7590 1910 7642
rect 1972 7590 1974 7642
rect 1812 7588 1836 7590
rect 1892 7588 1916 7590
rect 1972 7588 1996 7590
rect 1756 7568 2052 7588
rect 4756 7644 5052 7664
rect 4812 7642 4836 7644
rect 4892 7642 4916 7644
rect 4972 7642 4996 7644
rect 4834 7590 4836 7642
rect 4898 7590 4910 7642
rect 4972 7590 4974 7642
rect 4812 7588 4836 7590
rect 4892 7588 4916 7590
rect 4972 7588 4996 7590
rect 4756 7568 5052 7588
rect 6104 7342 6132 8230
rect 6196 7886 6224 8774
rect 6256 8188 6552 8208
rect 6312 8186 6336 8188
rect 6392 8186 6416 8188
rect 6472 8186 6496 8188
rect 6334 8134 6336 8186
rect 6398 8134 6410 8186
rect 6472 8134 6474 8186
rect 6312 8132 6336 8134
rect 6392 8132 6416 8134
rect 6472 8132 6496 8134
rect 6256 8112 6552 8132
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 3256 7100 3552 7120
rect 3312 7098 3336 7100
rect 3392 7098 3416 7100
rect 3472 7098 3496 7100
rect 3334 7046 3336 7098
rect 3398 7046 3410 7098
rect 3472 7046 3474 7098
rect 3312 7044 3336 7046
rect 3392 7044 3416 7046
rect 3472 7044 3496 7046
rect 3256 7024 3552 7044
rect 6104 6780 6132 7278
rect 6256 7100 6552 7120
rect 6312 7098 6336 7100
rect 6392 7098 6416 7100
rect 6472 7098 6496 7100
rect 6334 7046 6336 7098
rect 6398 7046 6410 7098
rect 6472 7046 6474 7098
rect 6312 7044 6336 7046
rect 6392 7044 6416 7046
rect 6472 7044 6496 7046
rect 6256 7024 6552 7044
rect 6276 6792 6328 6798
rect 6104 6752 6276 6780
rect 6276 6734 6328 6740
rect 1756 6556 2052 6576
rect 1812 6554 1836 6556
rect 1892 6554 1916 6556
rect 1972 6554 1996 6556
rect 1834 6502 1836 6554
rect 1898 6502 1910 6554
rect 1972 6502 1974 6554
rect 1812 6500 1836 6502
rect 1892 6500 1916 6502
rect 1972 6500 1996 6502
rect 1756 6480 2052 6500
rect 4756 6556 5052 6576
rect 4812 6554 4836 6556
rect 4892 6554 4916 6556
rect 4972 6554 4996 6556
rect 4834 6502 4836 6554
rect 4898 6502 4910 6554
rect 4972 6502 4974 6554
rect 4812 6500 4836 6502
rect 4892 6500 4916 6502
rect 4972 6500 4996 6502
rect 4756 6480 5052 6500
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 3256 6012 3552 6032
rect 3312 6010 3336 6012
rect 3392 6010 3416 6012
rect 3472 6010 3496 6012
rect 3334 5958 3336 6010
rect 3398 5958 3410 6010
rect 3472 5958 3474 6010
rect 3312 5956 3336 5958
rect 3392 5956 3416 5958
rect 3472 5956 3496 5958
rect 3256 5936 3552 5956
rect 5368 5914 5396 6326
rect 6288 6322 6316 6734
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 5552 5914 5580 6258
rect 6256 6012 6552 6032
rect 6312 6010 6336 6012
rect 6392 6010 6416 6012
rect 6472 6010 6496 6012
rect 6334 5958 6336 6010
rect 6398 5958 6410 6010
rect 6472 5958 6474 6010
rect 6312 5956 6336 5958
rect 6392 5956 6416 5958
rect 6472 5956 6496 5958
rect 6256 5936 6552 5956
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6656 5642 6684 6598
rect 6748 5778 6776 8978
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7116 8090 7144 8366
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7546 7052 7822
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7116 7478 7144 8026
rect 7392 7546 7420 8570
rect 7576 8362 7604 9590
rect 7668 8566 7696 10406
rect 7756 9820 8052 9840
rect 7812 9818 7836 9820
rect 7892 9818 7916 9820
rect 7972 9818 7996 9820
rect 7834 9766 7836 9818
rect 7898 9766 7910 9818
rect 7972 9766 7974 9818
rect 7812 9764 7836 9766
rect 7892 9764 7916 9766
rect 7972 9764 7996 9766
rect 7756 9744 8052 9764
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7760 9110 7788 9590
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 8128 8974 8156 10746
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 10470 8340 10542
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10198 8340 10406
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9722 8340 9998
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8312 9178 8340 9658
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7756 8732 8052 8752
rect 7812 8730 7836 8732
rect 7892 8730 7916 8732
rect 7972 8730 7996 8732
rect 7834 8678 7836 8730
rect 7898 8678 7910 8730
rect 7972 8678 7974 8730
rect 7812 8676 7836 8678
rect 7892 8676 7916 8678
rect 7972 8676 7996 8678
rect 7756 8656 8052 8676
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 8312 7954 8340 8434
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 7472 7812 7524 7818
rect 7472 7754 7524 7760
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7484 6798 7512 7754
rect 7756 7644 8052 7664
rect 7812 7642 7836 7644
rect 7892 7642 7916 7644
rect 7972 7642 7996 7644
rect 7834 7590 7836 7642
rect 7898 7590 7910 7642
rect 7972 7590 7974 7642
rect 7812 7588 7836 7590
rect 7892 7588 7916 7590
rect 7972 7588 7996 7590
rect 7756 7568 8052 7588
rect 8312 7546 8340 7890
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6840 5914 6868 6666
rect 7484 6458 7512 6734
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7668 6322 7696 6734
rect 7756 6556 8052 6576
rect 7812 6554 7836 6556
rect 7892 6554 7916 6556
rect 7972 6554 7996 6556
rect 7834 6502 7836 6554
rect 7898 6502 7910 6554
rect 7972 6502 7974 6554
rect 7812 6500 7836 6502
rect 7892 6500 7916 6502
rect 7972 6500 7996 6502
rect 7756 6480 8052 6500
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8300 6316 8352 6322
rect 8404 6304 8432 12378
rect 11060 12300 11112 12306
rect 11112 12260 11192 12288
rect 11060 12242 11112 12248
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11898 10640 12038
rect 10756 11996 11052 12016
rect 10812 11994 10836 11996
rect 10892 11994 10916 11996
rect 10972 11994 10996 11996
rect 10834 11942 10836 11994
rect 10898 11942 10910 11994
rect 10972 11942 10974 11994
rect 10812 11940 10836 11942
rect 10892 11940 10916 11942
rect 10972 11940 10996 11942
rect 10756 11920 11052 11940
rect 11164 11898 11192 12260
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8956 11014 8984 11698
rect 9256 11452 9552 11472
rect 9312 11450 9336 11452
rect 9392 11450 9416 11452
rect 9472 11450 9496 11452
rect 9334 11398 9336 11450
rect 9398 11398 9410 11450
rect 9472 11398 9474 11450
rect 9312 11396 9336 11398
rect 9392 11396 9416 11398
rect 9472 11396 9496 11398
rect 9256 11376 9552 11396
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10674 8984 10950
rect 9048 10674 9076 11086
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 9048 10266 9076 10610
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 8566 8616 9998
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8680 9042 8708 9658
rect 9140 9450 9168 10474
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9256 10364 9552 10384
rect 9312 10362 9336 10364
rect 9392 10362 9416 10364
rect 9472 10362 9496 10364
rect 9334 10310 9336 10362
rect 9398 10310 9410 10362
rect 9472 10310 9474 10362
rect 9312 10308 9336 10310
rect 9392 10308 9416 10310
rect 9472 10308 9496 10310
rect 9256 10288 9552 10308
rect 9600 9518 9628 10406
rect 10336 9926 10364 10610
rect 10428 10130 10456 11766
rect 10612 10248 10640 11834
rect 11256 11694 11284 12922
rect 11900 12306 11928 13942
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12256 13628 12552 13648
rect 12312 13626 12336 13628
rect 12392 13626 12416 13628
rect 12472 13626 12496 13628
rect 12334 13574 12336 13626
rect 12398 13574 12410 13626
rect 12472 13574 12474 13626
rect 12312 13572 12336 13574
rect 12392 13572 12416 13574
rect 12472 13572 12496 13574
rect 12256 13552 12552 13572
rect 12728 13190 12756 13738
rect 12912 13530 12940 14282
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 13096 13394 13124 13874
rect 13280 13462 13308 13874
rect 13464 13802 13492 13874
rect 13452 13796 13504 13802
rect 13648 13784 13676 14758
rect 13832 14346 13860 14962
rect 14200 14482 14228 15302
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14618 14596 14962
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14660 14550 14688 15302
rect 15396 15162 15424 15438
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15488 15094 15516 15370
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 14648 14544 14700 14550
rect 14648 14486 14700 14492
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 13756 14172 14052 14192
rect 13812 14170 13836 14172
rect 13892 14170 13916 14172
rect 13972 14170 13996 14172
rect 13834 14118 13836 14170
rect 13898 14118 13910 14170
rect 13972 14118 13974 14170
rect 13812 14116 13836 14118
rect 13892 14116 13916 14118
rect 13972 14116 13996 14118
rect 13756 14096 14052 14116
rect 14292 13870 14320 14282
rect 14844 13938 14872 15030
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15028 14006 15056 14962
rect 15256 14716 15552 14736
rect 15312 14714 15336 14716
rect 15392 14714 15416 14716
rect 15472 14714 15496 14716
rect 15334 14662 15336 14714
rect 15398 14662 15410 14714
rect 15472 14662 15474 14714
rect 15312 14660 15336 14662
rect 15392 14660 15416 14662
rect 15472 14660 15496 14662
rect 15256 14640 15552 14660
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15016 14000 15068 14006
rect 15016 13942 15068 13948
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 13728 13796 13780 13802
rect 13648 13756 13728 13784
rect 13452 13738 13504 13744
rect 13728 13738 13780 13744
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13740 13326 13768 13738
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 13452 13320 13504 13326
rect 13728 13320 13780 13326
rect 13452 13262 13504 13268
rect 13648 13280 13728 13308
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12256 12540 12552 12560
rect 12312 12538 12336 12540
rect 12392 12538 12416 12540
rect 12472 12538 12496 12540
rect 12334 12486 12336 12538
rect 12398 12486 12410 12538
rect 12472 12486 12474 12538
rect 12312 12484 12336 12486
rect 12392 12484 12416 12486
rect 12472 12484 12496 12486
rect 12256 12464 12552 12484
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11348 11898 11376 12106
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11808 11830 11836 12106
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11808 11354 11836 11766
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10756 10908 11052 10928
rect 10812 10906 10836 10908
rect 10892 10906 10916 10908
rect 10972 10906 10996 10908
rect 10834 10854 10836 10906
rect 10898 10854 10910 10906
rect 10972 10854 10974 10906
rect 10812 10852 10836 10854
rect 10892 10852 10916 10854
rect 10972 10852 10996 10854
rect 10756 10832 11052 10852
rect 11164 10810 11192 11086
rect 11152 10804 11204 10810
rect 11204 10764 11284 10792
rect 11152 10746 11204 10752
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10692 10260 10744 10266
rect 10612 10220 10692 10248
rect 10692 10202 10744 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9140 9178 9168 9386
rect 9256 9276 9552 9296
rect 9312 9274 9336 9276
rect 9392 9274 9416 9276
rect 9472 9274 9496 9276
rect 9334 9222 9336 9274
rect 9398 9222 9410 9274
rect 9472 9222 9474 9274
rect 9312 9220 9336 9222
rect 9392 9220 9416 9222
rect 9472 9220 9496 9222
rect 9256 9200 9552 9220
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8772 8022 8800 8570
rect 9600 8430 9628 9454
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9048 8090 9076 8366
rect 9256 8188 9552 8208
rect 9312 8186 9336 8188
rect 9392 8186 9416 8188
rect 9472 8186 9496 8188
rect 9334 8134 9336 8186
rect 9398 8134 9410 8186
rect 9472 8134 9474 8186
rect 9312 8132 9336 8134
rect 9392 8132 9416 8134
rect 9472 8132 9496 8134
rect 9256 8112 9552 8132
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8772 7886 8800 7958
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 9140 7410 9168 8026
rect 9600 7886 9628 8366
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9876 7546 9904 8842
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9140 6934 9168 7346
rect 9256 7100 9552 7120
rect 9312 7098 9336 7100
rect 9392 7098 9416 7100
rect 9472 7098 9496 7100
rect 9334 7046 9336 7098
rect 9398 7046 9410 7098
rect 9472 7046 9474 7098
rect 9312 7044 9336 7046
rect 9392 7044 9416 7046
rect 9472 7044 9496 7046
rect 9256 7024 9552 7044
rect 9876 7002 9904 7482
rect 9968 7478 9996 7822
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10060 7206 10088 8502
rect 10152 8022 10180 8910
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8090 10272 8842
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 7886 10180 7958
rect 10336 7886 10364 9862
rect 10428 9722 10456 10066
rect 11164 9994 11192 10474
rect 10600 9988 10652 9994
rect 10600 9930 10652 9936
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9042 10548 9522
rect 10612 9518 10640 9930
rect 10756 9820 11052 9840
rect 10812 9818 10836 9820
rect 10892 9818 10916 9820
rect 10972 9818 10996 9820
rect 10834 9766 10836 9818
rect 10898 9766 10910 9818
rect 10972 9766 10974 9818
rect 10812 9764 10836 9766
rect 10892 9764 10916 9766
rect 10972 9764 10996 9766
rect 10756 9744 11052 9764
rect 11164 9722 11192 9930
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11256 9654 11284 10764
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 11152 9512 11204 9518
rect 11348 9500 11376 11154
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10810 11652 10950
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11900 10674 11928 12242
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12256 11452 12552 11472
rect 12312 11450 12336 11452
rect 12392 11450 12416 11452
rect 12472 11450 12496 11452
rect 12334 11398 12336 11450
rect 12398 11398 12410 11450
rect 12472 11398 12474 11450
rect 12312 11396 12336 11398
rect 12392 11396 12416 11398
rect 12472 11396 12496 11398
rect 12256 11376 12552 11396
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11992 10470 12020 11086
rect 12636 10742 12664 11630
rect 12728 11218 12756 13126
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 11762 13216 12242
rect 13280 12238 13308 12786
rect 13464 12782 13492 13262
rect 13648 12986 13676 13280
rect 13728 13262 13780 13268
rect 13756 13084 14052 13104
rect 13812 13082 13836 13084
rect 13892 13082 13916 13084
rect 13972 13082 13996 13084
rect 13834 13030 13836 13082
rect 13898 13030 13910 13082
rect 13972 13030 13974 13082
rect 13812 13028 13836 13030
rect 13892 13028 13916 13030
rect 13972 13028 13996 13030
rect 13756 13008 14052 13028
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 14200 12918 14228 13330
rect 14292 13326 14320 13806
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13464 12102 13492 12718
rect 13556 12714 13584 12786
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13556 12442 13584 12650
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13188 11354 13216 11698
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13464 11218 13492 11698
rect 13556 11694 13584 12106
rect 13756 11996 14052 12016
rect 13812 11994 13836 11996
rect 13892 11994 13916 11996
rect 13972 11994 13996 11996
rect 13834 11942 13836 11994
rect 13898 11942 13910 11994
rect 13972 11942 13974 11994
rect 13812 11940 13836 11942
rect 13892 11940 13916 11942
rect 13972 11940 13996 11942
rect 13756 11920 14052 11940
rect 14108 11762 14136 12718
rect 14292 12288 14320 13262
rect 14752 13258 14780 13874
rect 14844 13530 14872 13874
rect 15028 13530 15056 13942
rect 15120 13938 15148 14554
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 15120 13462 15148 13874
rect 15256 13628 15552 13648
rect 15312 13626 15336 13628
rect 15392 13626 15416 13628
rect 15472 13626 15496 13628
rect 15334 13574 15336 13626
rect 15398 13574 15410 13626
rect 15472 13574 15474 13626
rect 15312 13572 15336 13574
rect 15392 13572 15416 13574
rect 15472 13572 15496 13574
rect 15256 13552 15552 13572
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14200 12260 14320 12288
rect 14200 11830 14228 12260
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13556 10810 13584 11630
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11286 13768 11562
rect 14108 11354 14136 11698
rect 14292 11694 14320 12106
rect 14476 11898 14504 12174
rect 14660 12102 14688 12718
rect 14752 12322 14780 13194
rect 14752 12294 14872 12322
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 13728 11280 13780 11286
rect 13648 11240 13728 11268
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 11992 10198 12020 10406
rect 12256 10364 12552 10384
rect 12312 10362 12336 10364
rect 12392 10362 12416 10364
rect 12472 10362 12496 10364
rect 12334 10310 12336 10362
rect 12398 10310 12410 10362
rect 12472 10310 12474 10362
rect 12312 10308 12336 10310
rect 12392 10308 12416 10310
rect 12472 10308 12496 10310
rect 12256 10288 12552 10308
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11900 9586 11928 9658
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11204 9472 11376 9500
rect 11152 9454 11204 9460
rect 10612 9178 10640 9454
rect 10796 9178 10824 9454
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10756 8732 11052 8752
rect 10812 8730 10836 8732
rect 10892 8730 10916 8732
rect 10972 8730 10996 8732
rect 10834 8678 10836 8730
rect 10898 8678 10910 8730
rect 10972 8678 10974 8730
rect 10812 8676 10836 8678
rect 10892 8676 10916 8678
rect 10972 8676 10996 8678
rect 10756 8656 11052 8676
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 7954 10824 8366
rect 11164 8362 11192 9454
rect 11532 8634 11560 9522
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11808 8634 11836 8842
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10152 7478 10180 7822
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 10244 7546 10272 7754
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10336 7342 10364 7822
rect 10756 7644 11052 7664
rect 10812 7642 10836 7644
rect 10892 7642 10916 7644
rect 10972 7642 10996 7644
rect 10834 7590 10836 7642
rect 10898 7590 10910 7642
rect 10972 7590 10974 7642
rect 10812 7588 10836 7590
rect 10892 7588 10916 7590
rect 10972 7588 10996 7590
rect 10756 7568 11052 7588
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 8352 6276 8432 6304
rect 8760 6316 8812 6322
rect 8300 6258 8352 6264
rect 8760 6258 8812 6264
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 1756 5468 2052 5488
rect 1812 5466 1836 5468
rect 1892 5466 1916 5468
rect 1972 5466 1996 5468
rect 1834 5414 1836 5466
rect 1898 5414 1910 5466
rect 1972 5414 1974 5466
rect 1812 5412 1836 5414
rect 1892 5412 1916 5414
rect 1972 5412 1996 5414
rect 1756 5392 2052 5412
rect 4756 5468 5052 5488
rect 4812 5466 4836 5468
rect 4892 5466 4916 5468
rect 4972 5466 4996 5468
rect 4834 5414 4836 5466
rect 4898 5414 4910 5466
rect 4972 5414 4974 5466
rect 4812 5412 4836 5414
rect 4892 5412 4916 5414
rect 4972 5412 4996 5414
rect 4756 5392 5052 5412
rect 6656 5370 6684 5578
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6748 5234 6776 5714
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 3256 4924 3552 4944
rect 3312 4922 3336 4924
rect 3392 4922 3416 4924
rect 3472 4922 3496 4924
rect 3334 4870 3336 4922
rect 3398 4870 3410 4922
rect 3472 4870 3474 4922
rect 3312 4868 3336 4870
rect 3392 4868 3416 4870
rect 3472 4868 3496 4870
rect 3256 4848 3552 4868
rect 6256 4924 6552 4944
rect 6312 4922 6336 4924
rect 6392 4922 6416 4924
rect 6472 4922 6496 4924
rect 6334 4870 6336 4922
rect 6398 4870 6410 4922
rect 6472 4870 6474 4922
rect 6312 4868 6336 4870
rect 6392 4868 6416 4870
rect 6472 4868 6496 4870
rect 6256 4848 6552 4868
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 1756 4380 2052 4400
rect 1812 4378 1836 4380
rect 1892 4378 1916 4380
rect 1972 4378 1996 4380
rect 1834 4326 1836 4378
rect 1898 4326 1910 4378
rect 1972 4326 1974 4378
rect 1812 4324 1836 4326
rect 1892 4324 1916 4326
rect 1972 4324 1996 4326
rect 1756 4304 2052 4324
rect 4756 4380 5052 4400
rect 4812 4378 4836 4380
rect 4892 4378 4916 4380
rect 4972 4378 4996 4380
rect 4834 4326 4836 4378
rect 4898 4326 4910 4378
rect 4972 4326 4974 4378
rect 4812 4324 4836 4326
rect 4892 4324 4916 4326
rect 4972 4324 4996 4326
rect 4756 4304 5052 4324
rect 6656 3942 6684 4422
rect 6748 4214 6776 5170
rect 6840 4826 6868 5850
rect 7024 5778 7052 6190
rect 7668 5914 7696 6258
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7024 5370 7052 5714
rect 7756 5468 8052 5488
rect 7812 5466 7836 5468
rect 7892 5466 7916 5468
rect 7972 5466 7996 5468
rect 7834 5414 7836 5466
rect 7898 5414 7910 5466
rect 7972 5414 7974 5466
rect 7812 5412 7836 5414
rect 7892 5412 7916 5414
rect 7972 5412 7996 5414
rect 7756 5392 8052 5412
rect 8128 5370 8156 6258
rect 8312 6186 8340 6258
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8312 5302 8340 6122
rect 8680 5574 8708 6190
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5302 8708 5510
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8772 4826 8800 6258
rect 9140 5778 9168 6870
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9256 6012 9552 6032
rect 9312 6010 9336 6012
rect 9392 6010 9416 6012
rect 9472 6010 9496 6012
rect 9334 5958 9336 6010
rect 9398 5958 9410 6010
rect 9472 5958 9474 6010
rect 9312 5956 9336 5958
rect 9392 5956 9416 5958
rect 9472 5956 9496 5958
rect 9256 5936 9552 5956
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9140 5302 9168 5714
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9600 5234 9628 6394
rect 9876 6390 9904 6938
rect 10060 6798 10088 7142
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6458 10088 6734
rect 10612 6458 10640 7142
rect 10888 7002 10916 7278
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10756 6556 11052 6576
rect 10812 6554 10836 6556
rect 10892 6554 10916 6556
rect 10972 6554 10996 6556
rect 10834 6502 10836 6554
rect 10898 6502 10910 6554
rect 10972 6502 10974 6554
rect 10812 6500 10836 6502
rect 10892 6500 10916 6502
rect 10972 6500 10996 6502
rect 10756 6480 11052 6500
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9968 5710 9996 6258
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9140 4826 9168 5034
rect 9256 4924 9552 4944
rect 9312 4922 9336 4924
rect 9392 4922 9416 4924
rect 9472 4922 9496 4924
rect 9334 4870 9336 4922
rect 9398 4870 9410 4922
rect 9472 4870 9474 4922
rect 9312 4868 9336 4870
rect 9392 4868 9416 4870
rect 9472 4868 9496 4870
rect 9256 4848 9552 4868
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9600 4622 9628 5170
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 7756 4380 8052 4400
rect 7812 4378 7836 4380
rect 7892 4378 7916 4380
rect 7972 4378 7996 4380
rect 7834 4326 7836 4378
rect 7898 4326 7910 4378
rect 7972 4326 7974 4378
rect 7812 4324 7836 4326
rect 7892 4324 7916 4326
rect 7972 4324 7996 4326
rect 7756 4304 8052 4324
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 8128 4154 8156 4490
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 8036 4126 8156 4154
rect 7668 4049 7696 4082
rect 7654 4040 7710 4049
rect 7654 3975 7710 3984
rect 8036 3942 8064 4126
rect 8312 3942 8340 4558
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 3256 3836 3552 3856
rect 3312 3834 3336 3836
rect 3392 3834 3416 3836
rect 3472 3834 3496 3836
rect 3334 3782 3336 3834
rect 3398 3782 3410 3834
rect 3472 3782 3474 3834
rect 3312 3780 3336 3782
rect 3392 3780 3416 3782
rect 3472 3780 3496 3782
rect 3256 3760 3552 3780
rect 6256 3836 6552 3856
rect 6312 3834 6336 3836
rect 6392 3834 6416 3836
rect 6472 3834 6496 3836
rect 6334 3782 6336 3834
rect 6398 3782 6410 3834
rect 6472 3782 6474 3834
rect 6312 3780 6336 3782
rect 6392 3780 6416 3782
rect 6472 3780 6496 3782
rect 6256 3760 6552 3780
rect 1756 3292 2052 3312
rect 1812 3290 1836 3292
rect 1892 3290 1916 3292
rect 1972 3290 1996 3292
rect 1834 3238 1836 3290
rect 1898 3238 1910 3290
rect 1972 3238 1974 3290
rect 1812 3236 1836 3238
rect 1892 3236 1916 3238
rect 1972 3236 1996 3238
rect 1756 3216 2052 3236
rect 4756 3292 5052 3312
rect 4812 3290 4836 3292
rect 4892 3290 4916 3292
rect 4972 3290 4996 3292
rect 4834 3238 4836 3290
rect 4898 3238 4910 3290
rect 4972 3238 4974 3290
rect 4812 3236 4836 3238
rect 4892 3236 4916 3238
rect 4972 3236 4996 3238
rect 4756 3216 5052 3236
rect 6656 3194 6684 3878
rect 7208 3738 7236 3878
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 8036 3670 8064 3878
rect 8024 3664 8076 3670
rect 8076 3624 8156 3652
rect 8024 3606 8076 3612
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 7392 3058 7420 3334
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 3256 2748 3552 2768
rect 3312 2746 3336 2748
rect 3392 2746 3416 2748
rect 3472 2746 3496 2748
rect 3334 2694 3336 2746
rect 3398 2694 3410 2746
rect 3472 2694 3474 2746
rect 3312 2692 3336 2694
rect 3392 2692 3416 2694
rect 3472 2692 3496 2694
rect 3256 2672 3552 2692
rect 6256 2748 6552 2768
rect 6312 2746 6336 2748
rect 6392 2746 6416 2748
rect 6472 2746 6496 2748
rect 6334 2694 6336 2746
rect 6398 2694 6410 2746
rect 6472 2694 6474 2746
rect 6312 2692 6336 2694
rect 6392 2692 6416 2694
rect 6472 2692 6496 2694
rect 6256 2672 6552 2692
rect 7300 2446 7328 2994
rect 7668 2650 7696 3538
rect 7756 3292 8052 3312
rect 7812 3290 7836 3292
rect 7892 3290 7916 3292
rect 7972 3290 7996 3292
rect 7834 3238 7836 3290
rect 7898 3238 7910 3290
rect 7972 3238 7974 3290
rect 7812 3236 7836 3238
rect 7892 3236 7916 3238
rect 7972 3236 7996 3238
rect 7756 3216 8052 3236
rect 8128 3194 8156 3624
rect 8312 3534 8340 3878
rect 8496 3602 8524 4422
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8484 3460 8536 3466
rect 8588 3448 8616 4014
rect 8536 3420 8616 3448
rect 8484 3402 8536 3408
rect 8588 3194 8616 3420
rect 8864 3398 8892 4150
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 9048 3194 9076 4150
rect 9508 3924 9536 4490
rect 9588 3936 9640 3942
rect 9508 3896 9588 3924
rect 9588 3878 9640 3884
rect 9256 3836 9552 3856
rect 9312 3834 9336 3836
rect 9392 3834 9416 3836
rect 9472 3834 9496 3836
rect 9334 3782 9336 3834
rect 9398 3782 9410 3834
rect 9472 3782 9474 3834
rect 9312 3780 9336 3782
rect 9392 3780 9416 3782
rect 9472 3780 9496 3782
rect 9256 3760 9552 3780
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 9140 2378 9168 2994
rect 9508 2990 9536 3334
rect 9784 3126 9812 3402
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9496 2984 9548 2990
rect 9548 2944 9628 2972
rect 9496 2926 9548 2932
rect 9256 2748 9552 2768
rect 9312 2746 9336 2748
rect 9392 2746 9416 2748
rect 9472 2746 9496 2748
rect 9334 2694 9336 2746
rect 9398 2694 9410 2746
rect 9472 2694 9474 2746
rect 9312 2692 9336 2694
rect 9392 2692 9416 2694
rect 9472 2692 9496 2694
rect 9256 2672 9552 2692
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9600 2310 9628 2944
rect 9784 2650 9812 3062
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 1756 2204 2052 2224
rect 1812 2202 1836 2204
rect 1892 2202 1916 2204
rect 1972 2202 1996 2204
rect 1834 2150 1836 2202
rect 1898 2150 1910 2202
rect 1972 2150 1974 2202
rect 1812 2148 1836 2150
rect 1892 2148 1916 2150
rect 1972 2148 1996 2150
rect 1756 2128 2052 2148
rect 4756 2204 5052 2224
rect 4812 2202 4836 2204
rect 4892 2202 4916 2204
rect 4972 2202 4996 2204
rect 4834 2150 4836 2202
rect 4898 2150 4910 2202
rect 4972 2150 4974 2202
rect 4812 2148 4836 2150
rect 4892 2148 4916 2150
rect 4972 2148 4996 2150
rect 4756 2128 5052 2148
rect 7756 2204 8052 2224
rect 7812 2202 7836 2204
rect 7892 2202 7916 2204
rect 7972 2202 7996 2204
rect 7834 2150 7836 2202
rect 7898 2150 7910 2202
rect 7972 2150 7974 2202
rect 7812 2148 7836 2150
rect 7892 2148 7916 2150
rect 7972 2148 7996 2150
rect 7756 2128 8052 2148
rect 18 60 74 800
rect 18 8 20 60
rect 72 8 74 60
rect 18 0 74 8
rect 9218 82 9274 800
rect 9324 82 9352 2246
rect 9218 54 9352 82
rect 9968 66 9996 5646
rect 10756 5468 11052 5488
rect 10812 5466 10836 5468
rect 10892 5466 10916 5468
rect 10972 5466 10996 5468
rect 10834 5414 10836 5466
rect 10898 5414 10910 5466
rect 10972 5414 10974 5466
rect 10812 5412 10836 5414
rect 10892 5412 10916 5414
rect 10972 5412 10996 5414
rect 10756 5392 11052 5412
rect 11164 5234 11192 7142
rect 11256 5642 11284 8366
rect 11440 8022 11468 8434
rect 11992 8430 12020 10134
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12176 8974 12204 9930
rect 13372 9654 13400 9998
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13372 9382 13400 9590
rect 13556 9518 13584 10610
rect 13648 9722 13676 11240
rect 13728 11222 13780 11228
rect 13756 10908 14052 10928
rect 13812 10906 13836 10908
rect 13892 10906 13916 10908
rect 13972 10906 13996 10908
rect 13834 10854 13836 10906
rect 13898 10854 13910 10906
rect 13972 10854 13974 10906
rect 13812 10852 13836 10854
rect 13892 10852 13916 10854
rect 13972 10852 13996 10854
rect 13756 10832 14052 10852
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10130 13860 10406
rect 14568 10266 14596 10678
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 13756 9820 14052 9840
rect 13812 9818 13836 9820
rect 13892 9818 13916 9820
rect 13972 9818 13996 9820
rect 13834 9766 13836 9818
rect 13898 9766 13910 9818
rect 13972 9766 13974 9818
rect 13812 9764 13836 9766
rect 13892 9764 13916 9766
rect 13972 9764 13996 9766
rect 13756 9744 14052 9764
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 14200 9518 14228 9862
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 12256 9276 12552 9296
rect 12312 9274 12336 9276
rect 12392 9274 12416 9276
rect 12472 9274 12496 9276
rect 12334 9222 12336 9274
rect 12398 9222 12410 9274
rect 12472 9222 12474 9274
rect 12312 9220 12336 9222
rect 12392 9220 12416 9222
rect 12472 9220 12496 9222
rect 12256 9200 12552 9220
rect 13556 9160 13584 9454
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 13372 9132 13584 9160
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13188 8430 13216 8842
rect 13372 8634 13400 9132
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13360 8628 13412 8634
rect 13280 8588 13360 8616
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 12256 8188 12552 8208
rect 12312 8186 12336 8188
rect 12392 8186 12416 8188
rect 12472 8186 12496 8188
rect 12334 8134 12336 8186
rect 12398 8134 12410 8186
rect 12472 8134 12474 8186
rect 12312 8132 12336 8134
rect 12392 8132 12416 8134
rect 12472 8132 12496 8134
rect 12256 8112 12552 8132
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11532 7478 11560 7686
rect 12268 7478 12296 7686
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6390 11744 6666
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11808 6322 11836 6938
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11348 5914 11376 6258
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 4049 10088 4626
rect 10244 4214 10272 4966
rect 11164 4622 11192 5170
rect 11256 5098 11284 5578
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4486 11192 4558
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 10756 4380 11052 4400
rect 10812 4378 10836 4380
rect 10892 4378 10916 4380
rect 10972 4378 10996 4380
rect 10834 4326 10836 4378
rect 10898 4326 10910 4378
rect 10972 4326 10974 4378
rect 10812 4324 10836 4326
rect 10892 4324 10916 4326
rect 10972 4324 10996 4326
rect 10756 4304 11052 4324
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10046 4040 10102 4049
rect 10046 3975 10102 3984
rect 10756 3292 11052 3312
rect 10812 3290 10836 3292
rect 10892 3290 10916 3292
rect 10972 3290 10996 3292
rect 10834 3238 10836 3290
rect 10898 3238 10910 3290
rect 10972 3238 10974 3290
rect 10812 3236 10836 3238
rect 10892 3236 10916 3238
rect 10972 3236 10996 3238
rect 10756 3216 11052 3236
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10244 2650 10272 3062
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 10060 2446 10088 2479
rect 11164 2446 11192 4082
rect 11348 3670 11376 5850
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11440 5234 11468 5578
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11428 4616 11480 4622
rect 11532 4604 11560 5510
rect 11624 5302 11652 5578
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11900 4826 11928 5170
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11900 4622 11928 4762
rect 12084 4622 12112 7142
rect 12256 7100 12552 7120
rect 12312 7098 12336 7100
rect 12392 7098 12416 7100
rect 12472 7098 12496 7100
rect 12334 7046 12336 7098
rect 12398 7046 12410 7098
rect 12472 7046 12474 7098
rect 12312 7044 12336 7046
rect 12392 7044 12416 7046
rect 12472 7044 12496 7046
rect 12256 7024 12552 7044
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12176 6458 12204 6666
rect 12728 6458 12756 7754
rect 12912 7478 12940 8366
rect 13188 8090 13216 8366
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 13280 7410 13308 8588
rect 13360 8570 13412 8576
rect 13464 8090 13492 8978
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 7546 13400 7822
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 7002 13308 7346
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13464 6866 13492 8026
rect 13556 7954 13584 8910
rect 13756 8732 14052 8752
rect 13812 8730 13836 8732
rect 13892 8730 13916 8732
rect 13972 8730 13996 8732
rect 13834 8678 13836 8730
rect 13898 8678 13910 8730
rect 13972 8678 13974 8730
rect 13812 8676 13836 8678
rect 13892 8676 13916 8678
rect 13972 8676 13996 8678
rect 13756 8656 14052 8676
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13556 7410 13584 7890
rect 13648 7750 13676 8502
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13756 7644 14052 7664
rect 13812 7642 13836 7644
rect 13892 7642 13916 7644
rect 13972 7642 13996 7644
rect 13834 7590 13836 7642
rect 13898 7590 13910 7642
rect 13972 7590 13974 7642
rect 13812 7588 13836 7590
rect 13892 7588 13916 7590
rect 13972 7588 13996 7590
rect 13756 7568 14052 7588
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 13464 6322 13492 6802
rect 13756 6556 14052 6576
rect 13812 6554 13836 6556
rect 13892 6554 13916 6556
rect 13972 6554 13996 6556
rect 13834 6502 13836 6554
rect 13898 6502 13910 6554
rect 13972 6502 13974 6554
rect 13812 6500 13836 6502
rect 13892 6500 13916 6502
rect 13972 6500 13996 6502
rect 13756 6480 14052 6500
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 12256 6012 12552 6032
rect 12312 6010 12336 6012
rect 12392 6010 12416 6012
rect 12472 6010 12496 6012
rect 12334 5958 12336 6010
rect 12398 5958 12410 6010
rect 12472 5958 12474 6010
rect 12312 5956 12336 5958
rect 12392 5956 12416 5958
rect 12472 5956 12496 5958
rect 12256 5936 12552 5956
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 13004 5710 13032 5782
rect 13096 5778 13124 6258
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12808 5704 12860 5710
rect 12992 5704 13044 5710
rect 12860 5664 12940 5692
rect 12808 5646 12860 5652
rect 12912 5234 12940 5664
rect 12992 5646 13044 5652
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12256 4924 12552 4944
rect 12312 4922 12336 4924
rect 12392 4922 12416 4924
rect 12472 4922 12496 4924
rect 12334 4870 12336 4922
rect 12398 4870 12410 4922
rect 12472 4870 12474 4922
rect 12312 4868 12336 4870
rect 12392 4868 12416 4870
rect 12472 4868 12496 4870
rect 12256 4848 12552 4868
rect 11480 4576 11560 4604
rect 11888 4616 11940 4622
rect 11428 4558 11480 4564
rect 11888 4558 11940 4564
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 11900 4282 11928 4558
rect 12728 4554 12756 5102
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11808 3738 11836 4150
rect 12728 4078 12756 4490
rect 12912 4214 12940 5170
rect 13004 5166 13032 5646
rect 13556 5574 13584 6190
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4214 13032 4422
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12256 3836 12552 3856
rect 12312 3834 12336 3836
rect 12392 3834 12416 3836
rect 12472 3834 12496 3836
rect 12334 3782 12336 3834
rect 12398 3782 12410 3834
rect 12472 3782 12474 3834
rect 12312 3780 12336 3782
rect 12392 3780 12416 3782
rect 12472 3780 12496 3782
rect 12256 3760 12552 3780
rect 12912 3738 12940 4150
rect 13188 4010 13216 4558
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13176 4004 13228 4010
rect 13096 3964 13176 3992
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11440 3602 11468 3674
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11256 2650 11284 3470
rect 11440 3194 11468 3538
rect 12912 3534 12940 3674
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 12636 3126 12664 3334
rect 13096 3194 13124 3964
rect 13176 3946 13228 3952
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12256 2748 12552 2768
rect 12312 2746 12336 2748
rect 12392 2746 12416 2748
rect 12472 2746 12496 2748
rect 12334 2694 12336 2746
rect 12398 2694 12410 2746
rect 12472 2694 12474 2746
rect 12312 2692 12336 2694
rect 12392 2692 12416 2694
rect 12472 2692 12496 2694
rect 12256 2672 12552 2692
rect 12912 2650 12940 2926
rect 13280 2650 13308 3062
rect 13372 2650 13400 4490
rect 13556 4282 13584 5510
rect 13756 5468 14052 5488
rect 13812 5466 13836 5468
rect 13892 5466 13916 5468
rect 13972 5466 13996 5468
rect 13834 5414 13836 5466
rect 13898 5414 13910 5466
rect 13972 5414 13974 5466
rect 13812 5412 13836 5414
rect 13892 5412 13916 5414
rect 13972 5412 13996 5414
rect 13756 5392 14052 5412
rect 14200 4570 14228 9318
rect 14476 8838 14504 9522
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 8566 14504 8774
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7478 14596 8230
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14292 5710 14320 7210
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6322 14412 7142
rect 14568 7002 14596 7414
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14660 6882 14688 12038
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 10606 14780 11630
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 10266 14780 10542
rect 14844 10266 14872 12294
rect 14936 11558 14964 13330
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15028 12374 15056 12786
rect 15580 12714 15608 15914
rect 15672 15026 15700 15982
rect 15764 15638 15792 16458
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14936 9722 14964 11494
rect 15028 11218 15056 12310
rect 15120 11762 15148 12582
rect 15256 12540 15552 12560
rect 15312 12538 15336 12540
rect 15392 12538 15416 12540
rect 15472 12538 15496 12540
rect 15334 12486 15336 12538
rect 15398 12486 15410 12538
rect 15472 12486 15474 12538
rect 15312 12484 15336 12486
rect 15392 12484 15416 12486
rect 15472 12484 15496 12486
rect 15256 12464 15552 12484
rect 15580 11762 15608 12650
rect 15672 11830 15700 13194
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15120 11354 15148 11698
rect 15256 11452 15552 11472
rect 15312 11450 15336 11452
rect 15392 11450 15416 11452
rect 15472 11450 15496 11452
rect 15334 11398 15336 11450
rect 15398 11398 15410 11450
rect 15472 11398 15474 11450
rect 15312 11396 15336 11398
rect 15392 11396 15416 11398
rect 15472 11396 15496 11398
rect 15256 11376 15552 11396
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15488 10742 15516 11086
rect 15580 11082 15608 11698
rect 15672 11286 15700 11766
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15764 10452 15792 13670
rect 15856 12850 15884 13806
rect 15948 13734 15976 14350
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 12442 15884 12786
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15948 12238 15976 13466
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 16040 11898 16068 15370
rect 16224 14414 16252 15506
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16224 14074 16252 14350
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16408 14006 16436 15302
rect 16500 14414 16528 16458
rect 16756 16348 17052 16368
rect 16812 16346 16836 16348
rect 16892 16346 16916 16348
rect 16972 16346 16996 16348
rect 16834 16294 16836 16346
rect 16898 16294 16910 16346
rect 16972 16294 16974 16346
rect 16812 16292 16836 16294
rect 16892 16292 16916 16294
rect 16972 16292 16996 16294
rect 16756 16272 17052 16292
rect 19756 16348 20052 16368
rect 19812 16346 19836 16348
rect 19892 16346 19916 16348
rect 19972 16346 19996 16348
rect 19834 16294 19836 16346
rect 19898 16294 19910 16346
rect 19972 16294 19974 16346
rect 19812 16292 19836 16294
rect 19892 16292 19916 16294
rect 19972 16292 19996 16294
rect 19756 16272 20052 16292
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 16592 15638 16620 15846
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16592 15026 16620 15574
rect 17328 15502 17356 15846
rect 18256 15804 18552 15824
rect 18312 15802 18336 15804
rect 18392 15802 18416 15804
rect 18472 15802 18496 15804
rect 18334 15750 18336 15802
rect 18398 15750 18410 15802
rect 18472 15750 18474 15802
rect 18312 15748 18336 15750
rect 18392 15748 18416 15750
rect 18472 15748 18496 15750
rect 18256 15728 18552 15748
rect 21256 15804 21552 15824
rect 21312 15802 21336 15804
rect 21392 15802 21416 15804
rect 21472 15802 21496 15804
rect 21334 15750 21336 15802
rect 21398 15750 21410 15802
rect 21472 15750 21474 15802
rect 21312 15748 21336 15750
rect 21392 15748 21416 15750
rect 21472 15748 21496 15750
rect 21256 15728 21552 15748
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 16756 15260 17052 15280
rect 16812 15258 16836 15260
rect 16892 15258 16916 15260
rect 16972 15258 16996 15260
rect 16834 15206 16836 15258
rect 16898 15206 16910 15258
rect 16972 15206 16974 15258
rect 16812 15204 16836 15206
rect 16892 15204 16916 15206
rect 16972 15204 16996 15206
rect 16756 15184 17052 15204
rect 17328 15094 17356 15438
rect 17788 15162 17816 15438
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16592 14618 16620 14962
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 17512 14550 17540 15030
rect 18156 14822 18184 15438
rect 18524 15094 18552 15438
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18800 14958 18828 15302
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 10588 16160 11630
rect 16224 11082 16252 13194
rect 16500 12986 16528 14350
rect 16756 14172 17052 14192
rect 16812 14170 16836 14172
rect 16892 14170 16916 14172
rect 16972 14170 16996 14172
rect 16834 14118 16836 14170
rect 16898 14118 16910 14170
rect 16972 14118 16974 14170
rect 16812 14116 16836 14118
rect 16892 14116 16916 14118
rect 16972 14116 16996 14118
rect 16756 14096 17052 14116
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16592 12986 16620 13738
rect 16684 13394 16712 13874
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16500 12238 16528 12718
rect 16684 12374 16712 13330
rect 17052 13326 17080 13942
rect 17144 13734 17172 14350
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17972 14006 18000 14214
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 18156 13870 18184 14758
rect 18256 14716 18552 14736
rect 18312 14714 18336 14716
rect 18392 14714 18416 14716
rect 18472 14714 18496 14716
rect 18334 14662 18336 14714
rect 18398 14662 18410 14714
rect 18472 14662 18474 14714
rect 18312 14660 18336 14662
rect 18392 14660 18416 14662
rect 18472 14660 18496 14662
rect 18256 14640 18552 14660
rect 18800 14414 18828 14894
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17040 13320 17092 13326
rect 17092 13280 17172 13308
rect 17040 13262 17092 13268
rect 16756 13084 17052 13104
rect 16812 13082 16836 13084
rect 16892 13082 16916 13084
rect 16972 13082 16996 13084
rect 16834 13030 16836 13082
rect 16898 13030 16910 13082
rect 16972 13030 16974 13082
rect 16812 13028 16836 13030
rect 16892 13028 16916 13030
rect 16972 13028 16996 13030
rect 16756 13008 17052 13028
rect 17144 12986 17172 13280
rect 18156 13190 18184 13806
rect 18256 13628 18552 13648
rect 18312 13626 18336 13628
rect 18392 13626 18416 13628
rect 18472 13626 18496 13628
rect 18334 13574 18336 13626
rect 18398 13574 18410 13626
rect 18472 13574 18474 13626
rect 18312 13572 18336 13574
rect 18392 13572 18416 13574
rect 18472 13572 18496 13574
rect 18256 13552 18552 13572
rect 18892 13258 18920 15098
rect 19168 14074 19196 15302
rect 19756 15260 20052 15280
rect 19812 15258 19836 15260
rect 19892 15258 19916 15260
rect 19972 15258 19996 15260
rect 19834 15206 19836 15258
rect 19898 15206 19910 15258
rect 19972 15206 19974 15258
rect 19812 15204 19836 15206
rect 19892 15204 19916 15206
rect 19972 15204 19996 15206
rect 19756 15184 20052 15204
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19444 14414 19472 14826
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19260 14074 19288 14350
rect 20364 14278 20392 14894
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 19756 14172 20052 14192
rect 19812 14170 19836 14172
rect 19892 14170 19916 14172
rect 19972 14170 19996 14172
rect 19834 14118 19836 14170
rect 19898 14118 19910 14170
rect 19972 14118 19974 14170
rect 19812 14116 19836 14118
rect 19892 14116 19916 14118
rect 19972 14116 19996 14118
rect 19756 14096 20052 14116
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19168 13938 19196 14010
rect 19260 13938 19564 13954
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19260 13932 19576 13938
rect 19260 13926 19524 13932
rect 19076 13326 19104 13874
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 18880 13252 18932 13258
rect 18880 13194 18932 13200
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 18064 12646 18092 13126
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11694 16528 12174
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16212 10600 16264 10606
rect 16132 10560 16212 10588
rect 16212 10542 16264 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15844 10464 15896 10470
rect 15764 10424 15844 10452
rect 15844 10406 15896 10412
rect 15256 10364 15552 10384
rect 15312 10362 15336 10364
rect 15392 10362 15416 10364
rect 15472 10362 15496 10364
rect 15334 10310 15336 10362
rect 15398 10310 15410 10362
rect 15472 10310 15474 10362
rect 15312 10308 15336 10310
rect 15392 10308 15416 10310
rect 15472 10308 15496 10310
rect 15256 10288 15552 10308
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9722 15424 9862
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15256 9276 15552 9296
rect 15312 9274 15336 9276
rect 15392 9274 15416 9276
rect 15472 9274 15496 9276
rect 15334 9222 15336 9274
rect 15398 9222 15410 9274
rect 15472 9222 15474 9274
rect 15312 9220 15336 9222
rect 15392 9220 15416 9222
rect 15472 9220 15496 9222
rect 15256 9200 15552 9220
rect 15672 8566 15700 9998
rect 15856 9518 15884 10406
rect 16224 10130 16252 10542
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15856 9042 15884 9454
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15256 8188 15552 8208
rect 15312 8186 15336 8188
rect 15392 8186 15416 8188
rect 15472 8186 15496 8188
rect 15334 8134 15336 8186
rect 15398 8134 15410 8186
rect 15472 8134 15474 8186
rect 15312 8132 15336 8134
rect 15392 8132 15416 8134
rect 15472 8132 15496 8134
rect 15256 8112 15552 8132
rect 15856 8090 15884 8434
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14832 7404 14884 7410
rect 15292 7404 15344 7410
rect 14832 7346 14884 7352
rect 15120 7364 15292 7392
rect 14752 7002 14780 7346
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14660 6854 14780 6882
rect 14844 6866 14872 7346
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14292 4690 14320 5646
rect 14384 5166 14412 6258
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5778 14504 6054
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14476 4826 14504 5714
rect 14660 5574 14688 6258
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14660 5234 14688 5510
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 4826 14688 5170
rect 14752 5030 14780 6854
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14936 5302 14964 7210
rect 15120 6934 15148 7364
rect 15292 7346 15344 7352
rect 15256 7100 15552 7120
rect 15312 7098 15336 7100
rect 15392 7098 15416 7100
rect 15472 7098 15496 7100
rect 15334 7046 15336 7098
rect 15398 7046 15410 7098
rect 15472 7046 15474 7098
rect 15312 7044 15336 7046
rect 15392 7044 15416 7046
rect 15472 7044 15496 7046
rect 15256 7024 15552 7044
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15672 6390 15700 6802
rect 15856 6798 15884 8026
rect 16040 7954 16068 9930
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16132 9178 16160 9522
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16132 7410 16160 9114
rect 16224 8090 16252 10066
rect 16316 9654 16344 10542
rect 16684 10266 16712 12310
rect 16756 11996 17052 12016
rect 16812 11994 16836 11996
rect 16892 11994 16916 11996
rect 16972 11994 16996 11996
rect 16834 11942 16836 11994
rect 16898 11942 16910 11994
rect 16972 11942 16974 11994
rect 16812 11940 16836 11942
rect 16892 11940 16916 11942
rect 16972 11940 16996 11942
rect 16756 11920 17052 11940
rect 17236 11830 17264 12582
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17604 11898 17632 12174
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11150 17172 11630
rect 17236 11286 17264 11766
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 16756 10908 17052 10928
rect 16812 10906 16836 10908
rect 16892 10906 16916 10908
rect 16972 10906 16996 10908
rect 16834 10854 16836 10906
rect 16898 10854 16910 10906
rect 16972 10854 16974 10906
rect 16812 10852 16836 10854
rect 16892 10852 16916 10854
rect 16972 10852 16996 10854
rect 16756 10832 17052 10852
rect 17328 10742 17356 11086
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16684 9994 16712 10202
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16756 9820 17052 9840
rect 16812 9818 16836 9820
rect 16892 9818 16916 9820
rect 16972 9818 16996 9820
rect 16834 9766 16836 9818
rect 16898 9766 16910 9818
rect 16972 9766 16974 9818
rect 16812 9764 16836 9766
rect 16892 9764 16916 9766
rect 16972 9764 16996 9766
rect 16756 9744 17052 9764
rect 17512 9654 17540 11494
rect 17604 11218 17632 11834
rect 17788 11830 17816 12174
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 10810 17724 11086
rect 17788 10810 17816 11766
rect 18064 11694 18092 12582
rect 18156 12238 18184 13126
rect 18892 12850 18920 13194
rect 19076 12850 19104 13262
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18256 12540 18552 12560
rect 18312 12538 18336 12540
rect 18392 12538 18416 12540
rect 18472 12538 18496 12540
rect 18334 12486 18336 12538
rect 18398 12486 18410 12538
rect 18472 12486 18474 12538
rect 18312 12484 18336 12486
rect 18392 12484 18416 12486
rect 18472 12484 18496 12486
rect 18256 12464 18552 12484
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 11354 18092 11630
rect 18156 11558 18184 12174
rect 18418 11792 18474 11801
rect 18708 11762 18736 12650
rect 18800 12102 18828 12786
rect 19168 12782 19196 13262
rect 19260 12986 19288 13926
rect 19524 13874 19576 13880
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13394 19380 13806
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 20364 13326 20392 14214
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20456 13530 20484 13874
rect 20548 13802 20576 15438
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14346 20668 14894
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20640 14074 20668 14282
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20536 13796 20588 13802
rect 20536 13738 20588 13744
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 19708 13320 19760 13326
rect 19628 13280 19708 13308
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 18418 11727 18474 11736
rect 18696 11756 18748 11762
rect 18432 11694 18460 11727
rect 18748 11716 18828 11744
rect 18696 11698 18748 11704
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18256 11452 18552 11472
rect 18312 11450 18336 11452
rect 18392 11450 18416 11452
rect 18472 11450 18496 11452
rect 18334 11398 18336 11450
rect 18398 11398 18410 11450
rect 18472 11398 18474 11450
rect 18312 11396 18336 11398
rect 18392 11396 18416 11398
rect 18472 11396 18496 11398
rect 18256 11376 18552 11396
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18800 11286 18828 11716
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 18256 10364 18552 10384
rect 18312 10362 18336 10364
rect 18392 10362 18416 10364
rect 18472 10362 18496 10364
rect 18334 10310 18336 10362
rect 18398 10310 18410 10362
rect 18472 10310 18474 10362
rect 18312 10308 18336 10310
rect 18392 10308 18416 10310
rect 18472 10308 18496 10310
rect 18256 10288 18552 10308
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16592 9178 16620 9522
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 17144 9042 17172 9318
rect 18256 9276 18552 9296
rect 18312 9274 18336 9276
rect 18392 9274 18416 9276
rect 18472 9274 18496 9276
rect 18334 9222 18336 9274
rect 18398 9222 18410 9274
rect 18472 9222 18474 9274
rect 18312 9220 18336 9222
rect 18392 9220 18416 9222
rect 18472 9220 18496 9222
rect 18256 9200 18552 9220
rect 18708 9178 18736 9930
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8634 16712 8910
rect 16756 8732 17052 8752
rect 16812 8730 16836 8732
rect 16892 8730 16916 8732
rect 16972 8730 16996 8732
rect 16834 8678 16836 8730
rect 16898 8678 16910 8730
rect 16972 8678 16974 8730
rect 16812 8676 16836 8678
rect 16892 8676 16916 8678
rect 16972 8676 16996 8678
rect 16756 8656 17052 8676
rect 17144 8634 17172 8978
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17696 8634 17724 8842
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 16684 8362 16712 8570
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16316 7750 16344 8230
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16120 7404 16172 7410
rect 16172 7364 16252 7392
rect 16120 7346 16172 7352
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6458 15884 6734
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15948 6322 15976 6666
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15256 6012 15552 6032
rect 15312 6010 15336 6012
rect 15392 6010 15416 6012
rect 15472 6010 15496 6012
rect 15334 5958 15336 6010
rect 15398 5958 15410 6010
rect 15472 5958 15474 6010
rect 15312 5956 15336 5958
rect 15392 5956 15416 5958
rect 15472 5956 15496 5958
rect 15256 5936 15552 5956
rect 15948 5710 15976 6258
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 5370 15976 5646
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 15256 4924 15552 4944
rect 15312 4922 15336 4924
rect 15392 4922 15416 4924
rect 15472 4922 15496 4924
rect 15334 4870 15336 4922
rect 15398 4870 15410 4922
rect 15472 4870 15474 4922
rect 15312 4868 15336 4870
rect 15392 4868 15416 4870
rect 15472 4868 15496 4870
rect 15256 4848 15552 4868
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 16040 4690 16068 5578
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 14372 4616 14424 4622
rect 14200 4564 14372 4570
rect 14200 4558 14424 4564
rect 14200 4542 14412 4558
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13648 3126 13676 4422
rect 13756 4380 14052 4400
rect 13812 4378 13836 4380
rect 13892 4378 13916 4380
rect 13972 4378 13996 4380
rect 13834 4326 13836 4378
rect 13898 4326 13910 4378
rect 13972 4326 13974 4378
rect 13812 4324 13836 4326
rect 13892 4324 13916 4326
rect 13972 4324 13996 4326
rect 13756 4304 14052 4324
rect 14384 4146 14412 4542
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13756 3292 14052 3312
rect 13812 3290 13836 3292
rect 13892 3290 13916 3292
rect 13972 3290 13996 3292
rect 13834 3238 13836 3290
rect 13898 3238 13910 3290
rect 13972 3238 13974 3290
rect 13812 3236 13836 3238
rect 13892 3236 13916 3238
rect 13972 3236 13996 3238
rect 13756 3216 14052 3236
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13648 2582 13676 3062
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13832 2446 13860 2790
rect 14108 2446 14136 3674
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 2854 14228 3334
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14292 2310 14320 3538
rect 14384 2922 14412 4082
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14476 3670 14504 3946
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14384 2553 14412 2858
rect 14568 2582 14596 3878
rect 14936 3126 14964 4014
rect 15028 3126 15056 4626
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15764 3942 15792 4422
rect 16040 4282 16068 4626
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15256 3836 15552 3856
rect 15312 3834 15336 3836
rect 15392 3834 15416 3836
rect 15472 3834 15496 3836
rect 15334 3782 15336 3834
rect 15398 3782 15410 3834
rect 15472 3782 15474 3834
rect 15312 3780 15336 3782
rect 15392 3780 15416 3782
rect 15472 3780 15496 3782
rect 15256 3760 15552 3780
rect 15764 3534 15792 3878
rect 16132 3534 16160 7142
rect 16224 5778 16252 7364
rect 16316 7002 16344 7686
rect 16684 7546 16712 7822
rect 16756 7644 17052 7664
rect 16812 7642 16836 7644
rect 16892 7642 16916 7644
rect 16972 7642 16996 7644
rect 16834 7590 16836 7642
rect 16898 7590 16910 7642
rect 16972 7590 16974 7642
rect 16812 7588 16836 7590
rect 16892 7588 16916 7590
rect 16972 7588 16996 7590
rect 16756 7568 17052 7588
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16684 7002 16712 7482
rect 17696 7002 17724 8570
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17788 7546 17816 8434
rect 18256 8188 18552 8208
rect 18312 8186 18336 8188
rect 18392 8186 18416 8188
rect 18472 8186 18496 8188
rect 18334 8134 18336 8186
rect 18398 8134 18410 8186
rect 18472 8134 18474 8186
rect 18312 8132 18336 8134
rect 18392 8132 18416 8134
rect 18472 8132 18496 8134
rect 18256 8112 18552 8132
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18248 7546 18276 7822
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18256 7100 18552 7120
rect 18312 7098 18336 7100
rect 18392 7098 18416 7100
rect 18472 7098 18496 7100
rect 18334 7046 18336 7098
rect 18398 7046 18410 7098
rect 18472 7046 18474 7098
rect 18312 7044 18336 7046
rect 18392 7044 18416 7046
rect 18472 7044 18496 7046
rect 18256 7024 18552 7044
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16224 5234 16252 5714
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16500 5030 16528 5646
rect 16592 5574 16620 6190
rect 16684 6118 16712 6734
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 16756 6556 17052 6576
rect 16812 6554 16836 6556
rect 16892 6554 16916 6556
rect 16972 6554 16996 6556
rect 16834 6502 16836 6554
rect 16898 6502 16910 6554
rect 16972 6502 16974 6554
rect 16812 6500 16836 6502
rect 16892 6500 16916 6502
rect 16972 6500 16996 6502
rect 16756 6480 17052 6500
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15764 2990 15792 3470
rect 16132 3194 16160 3470
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 15256 2748 15552 2768
rect 15312 2746 15336 2748
rect 15392 2746 15416 2748
rect 15472 2746 15496 2748
rect 15334 2694 15336 2746
rect 15398 2694 15410 2746
rect 15472 2694 15474 2746
rect 15312 2692 15336 2694
rect 15392 2692 15416 2694
rect 15472 2692 15496 2694
rect 15256 2672 15552 2692
rect 14556 2576 14608 2582
rect 14370 2544 14426 2553
rect 14556 2518 14608 2524
rect 14370 2479 14426 2488
rect 16316 2446 16344 4218
rect 16592 4010 16620 5510
rect 16684 5302 16712 6054
rect 17144 5710 17172 6190
rect 17972 5846 18000 6598
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 16756 5468 17052 5488
rect 16812 5466 16836 5468
rect 16892 5466 16916 5468
rect 16972 5466 16996 5468
rect 16834 5414 16836 5466
rect 16898 5414 16910 5466
rect 16972 5414 16974 5466
rect 16812 5412 16836 5414
rect 16892 5412 16916 5414
rect 16972 5412 16996 5414
rect 16756 5392 17052 5412
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17788 4690 17816 5102
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 17132 4616 17184 4622
rect 17132 4558 17184 4564
rect 16756 4380 17052 4400
rect 16812 4378 16836 4380
rect 16892 4378 16916 4380
rect 16972 4378 16996 4380
rect 16834 4326 16836 4378
rect 16898 4326 16910 4378
rect 16972 4326 16974 4378
rect 16812 4324 16836 4326
rect 16892 4324 16916 4326
rect 16972 4324 16996 4326
rect 16756 4304 17052 4324
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16868 3670 16896 4150
rect 17144 4010 17172 4558
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 17512 3602 17540 4082
rect 17788 4078 17816 4626
rect 17972 4146 18000 5646
rect 18156 4690 18184 6734
rect 18256 6012 18552 6032
rect 18312 6010 18336 6012
rect 18392 6010 18416 6012
rect 18472 6010 18496 6012
rect 18334 5958 18336 6010
rect 18398 5958 18410 6010
rect 18472 5958 18474 6010
rect 18312 5956 18336 5958
rect 18392 5956 18416 5958
rect 18472 5956 18496 5958
rect 18256 5936 18552 5956
rect 18616 5710 18644 8570
rect 18708 7818 18736 9114
rect 18800 8634 18828 11222
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 9042 18920 10610
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18984 9518 19012 10542
rect 19076 9926 19104 12038
rect 19168 11014 19196 12174
rect 19352 11801 19380 12786
rect 19628 12714 19656 13280
rect 19708 13262 19760 13268
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 19756 13084 20052 13104
rect 19812 13082 19836 13084
rect 19892 13082 19916 13084
rect 19972 13082 19996 13084
rect 19834 13030 19836 13082
rect 19898 13030 19910 13082
rect 19972 13030 19974 13082
rect 19812 13028 19836 13030
rect 19892 13028 19916 13030
rect 19972 13028 19996 13030
rect 19756 13008 20052 13028
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 20180 12442 20208 12854
rect 20732 12646 20760 14758
rect 21192 14618 21220 15030
rect 21256 14716 21552 14736
rect 21312 14714 21336 14716
rect 21392 14714 21416 14716
rect 21472 14714 21496 14716
rect 21334 14662 21336 14714
rect 21398 14662 21410 14714
rect 21472 14662 21474 14714
rect 21312 14660 21336 14662
rect 21392 14660 21416 14662
rect 21472 14660 21496 14662
rect 21256 14640 21552 14660
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21192 13734 21220 14350
rect 21652 13814 21680 27338
rect 22756 27228 23052 27248
rect 22812 27226 22836 27228
rect 22892 27226 22916 27228
rect 22972 27226 22996 27228
rect 22834 27174 22836 27226
rect 22898 27174 22910 27226
rect 22972 27174 22974 27226
rect 22812 27172 22836 27174
rect 22892 27172 22916 27174
rect 22972 27172 22996 27174
rect 22756 27152 23052 27172
rect 23124 27130 23152 27406
rect 25756 27228 26052 27248
rect 25812 27226 25836 27228
rect 25892 27226 25916 27228
rect 25972 27226 25996 27228
rect 25834 27174 25836 27226
rect 25898 27174 25910 27226
rect 25972 27174 25974 27226
rect 25812 27172 25836 27174
rect 25892 27172 25916 27174
rect 25972 27172 25996 27174
rect 25756 27152 26052 27172
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 24256 26684 24552 26704
rect 24312 26682 24336 26684
rect 24392 26682 24416 26684
rect 24472 26682 24496 26684
rect 24334 26630 24336 26682
rect 24398 26630 24410 26682
rect 24472 26630 24474 26682
rect 24312 26628 24336 26630
rect 24392 26628 24416 26630
rect 24472 26628 24496 26630
rect 24256 26608 24552 26628
rect 27256 26684 27552 26704
rect 27312 26682 27336 26684
rect 27392 26682 27416 26684
rect 27472 26682 27496 26684
rect 27334 26630 27336 26682
rect 27398 26630 27410 26682
rect 27472 26630 27474 26682
rect 27312 26628 27336 26630
rect 27392 26628 27416 26630
rect 27472 26628 27496 26630
rect 27256 26608 27552 26628
rect 22756 26140 23052 26160
rect 22812 26138 22836 26140
rect 22892 26138 22916 26140
rect 22972 26138 22996 26140
rect 22834 26086 22836 26138
rect 22898 26086 22910 26138
rect 22972 26086 22974 26138
rect 22812 26084 22836 26086
rect 22892 26084 22916 26086
rect 22972 26084 22996 26086
rect 22756 26064 23052 26084
rect 25756 26140 26052 26160
rect 25812 26138 25836 26140
rect 25892 26138 25916 26140
rect 25972 26138 25996 26140
rect 25834 26086 25836 26138
rect 25898 26086 25910 26138
rect 25972 26086 25974 26138
rect 25812 26084 25836 26086
rect 25892 26084 25916 26086
rect 25972 26084 25996 26086
rect 25756 26064 26052 26084
rect 24256 25596 24552 25616
rect 24312 25594 24336 25596
rect 24392 25594 24416 25596
rect 24472 25594 24496 25596
rect 24334 25542 24336 25594
rect 24398 25542 24410 25594
rect 24472 25542 24474 25594
rect 24312 25540 24336 25542
rect 24392 25540 24416 25542
rect 24472 25540 24496 25542
rect 24256 25520 24552 25540
rect 27256 25596 27552 25616
rect 27312 25594 27336 25596
rect 27392 25594 27416 25596
rect 27472 25594 27496 25596
rect 27334 25542 27336 25594
rect 27398 25542 27410 25594
rect 27472 25542 27474 25594
rect 27312 25540 27336 25542
rect 27392 25540 27416 25542
rect 27472 25540 27496 25542
rect 27256 25520 27552 25540
rect 22756 25052 23052 25072
rect 22812 25050 22836 25052
rect 22892 25050 22916 25052
rect 22972 25050 22996 25052
rect 22834 24998 22836 25050
rect 22898 24998 22910 25050
rect 22972 24998 22974 25050
rect 22812 24996 22836 24998
rect 22892 24996 22916 24998
rect 22972 24996 22996 24998
rect 22756 24976 23052 24996
rect 25756 25052 26052 25072
rect 25812 25050 25836 25052
rect 25892 25050 25916 25052
rect 25972 25050 25996 25052
rect 25834 24998 25836 25050
rect 25898 24998 25910 25050
rect 25972 24998 25974 25050
rect 25812 24996 25836 24998
rect 25892 24996 25916 24998
rect 25972 24996 25996 24998
rect 25756 24976 26052 24996
rect 24256 24508 24552 24528
rect 24312 24506 24336 24508
rect 24392 24506 24416 24508
rect 24472 24506 24496 24508
rect 24334 24454 24336 24506
rect 24398 24454 24410 24506
rect 24472 24454 24474 24506
rect 24312 24452 24336 24454
rect 24392 24452 24416 24454
rect 24472 24452 24496 24454
rect 24256 24432 24552 24452
rect 27256 24508 27552 24528
rect 27312 24506 27336 24508
rect 27392 24506 27416 24508
rect 27472 24506 27496 24508
rect 27334 24454 27336 24506
rect 27398 24454 27410 24506
rect 27472 24454 27474 24506
rect 27312 24452 27336 24454
rect 27392 24452 27416 24454
rect 27472 24452 27496 24454
rect 27256 24432 27552 24452
rect 22756 23964 23052 23984
rect 22812 23962 22836 23964
rect 22892 23962 22916 23964
rect 22972 23962 22996 23964
rect 22834 23910 22836 23962
rect 22898 23910 22910 23962
rect 22972 23910 22974 23962
rect 22812 23908 22836 23910
rect 22892 23908 22916 23910
rect 22972 23908 22996 23910
rect 22756 23888 23052 23908
rect 25756 23964 26052 23984
rect 25812 23962 25836 23964
rect 25892 23962 25916 23964
rect 25972 23962 25996 23964
rect 25834 23910 25836 23962
rect 25898 23910 25910 23962
rect 25972 23910 25974 23962
rect 25812 23908 25836 23910
rect 25892 23908 25916 23910
rect 25972 23908 25996 23910
rect 25756 23888 26052 23908
rect 24256 23420 24552 23440
rect 24312 23418 24336 23420
rect 24392 23418 24416 23420
rect 24472 23418 24496 23420
rect 24334 23366 24336 23418
rect 24398 23366 24410 23418
rect 24472 23366 24474 23418
rect 24312 23364 24336 23366
rect 24392 23364 24416 23366
rect 24472 23364 24496 23366
rect 24256 23344 24552 23364
rect 27256 23420 27552 23440
rect 27312 23418 27336 23420
rect 27392 23418 27416 23420
rect 27472 23418 27496 23420
rect 27334 23366 27336 23418
rect 27398 23366 27410 23418
rect 27472 23366 27474 23418
rect 27312 23364 27336 23366
rect 27392 23364 27416 23366
rect 27472 23364 27496 23366
rect 27256 23344 27552 23364
rect 22756 22876 23052 22896
rect 22812 22874 22836 22876
rect 22892 22874 22916 22876
rect 22972 22874 22996 22876
rect 22834 22822 22836 22874
rect 22898 22822 22910 22874
rect 22972 22822 22974 22874
rect 22812 22820 22836 22822
rect 22892 22820 22916 22822
rect 22972 22820 22996 22822
rect 22756 22800 23052 22820
rect 25756 22876 26052 22896
rect 25812 22874 25836 22876
rect 25892 22874 25916 22876
rect 25972 22874 25996 22876
rect 25834 22822 25836 22874
rect 25898 22822 25910 22874
rect 25972 22822 25974 22874
rect 25812 22820 25836 22822
rect 25892 22820 25916 22822
rect 25972 22820 25996 22822
rect 25756 22800 26052 22820
rect 24256 22332 24552 22352
rect 24312 22330 24336 22332
rect 24392 22330 24416 22332
rect 24472 22330 24496 22332
rect 24334 22278 24336 22330
rect 24398 22278 24410 22330
rect 24472 22278 24474 22330
rect 24312 22276 24336 22278
rect 24392 22276 24416 22278
rect 24472 22276 24496 22278
rect 24256 22256 24552 22276
rect 27256 22332 27552 22352
rect 27312 22330 27336 22332
rect 27392 22330 27416 22332
rect 27472 22330 27496 22332
rect 27334 22278 27336 22330
rect 27398 22278 27410 22330
rect 27472 22278 27474 22330
rect 27312 22276 27336 22278
rect 27392 22276 27416 22278
rect 27472 22276 27496 22278
rect 27256 22256 27552 22276
rect 22756 21788 23052 21808
rect 22812 21786 22836 21788
rect 22892 21786 22916 21788
rect 22972 21786 22996 21788
rect 22834 21734 22836 21786
rect 22898 21734 22910 21786
rect 22972 21734 22974 21786
rect 22812 21732 22836 21734
rect 22892 21732 22916 21734
rect 22972 21732 22996 21734
rect 22756 21712 23052 21732
rect 25756 21788 26052 21808
rect 25812 21786 25836 21788
rect 25892 21786 25916 21788
rect 25972 21786 25996 21788
rect 25834 21734 25836 21786
rect 25898 21734 25910 21786
rect 25972 21734 25974 21786
rect 25812 21732 25836 21734
rect 25892 21732 25916 21734
rect 25972 21732 25996 21734
rect 25756 21712 26052 21732
rect 24256 21244 24552 21264
rect 24312 21242 24336 21244
rect 24392 21242 24416 21244
rect 24472 21242 24496 21244
rect 24334 21190 24336 21242
rect 24398 21190 24410 21242
rect 24472 21190 24474 21242
rect 24312 21188 24336 21190
rect 24392 21188 24416 21190
rect 24472 21188 24496 21190
rect 24256 21168 24552 21188
rect 27256 21244 27552 21264
rect 27312 21242 27336 21244
rect 27392 21242 27416 21244
rect 27472 21242 27496 21244
rect 27334 21190 27336 21242
rect 27398 21190 27410 21242
rect 27472 21190 27474 21242
rect 27312 21188 27336 21190
rect 27392 21188 27416 21190
rect 27472 21188 27496 21190
rect 27256 21168 27552 21188
rect 22756 20700 23052 20720
rect 22812 20698 22836 20700
rect 22892 20698 22916 20700
rect 22972 20698 22996 20700
rect 22834 20646 22836 20698
rect 22898 20646 22910 20698
rect 22972 20646 22974 20698
rect 22812 20644 22836 20646
rect 22892 20644 22916 20646
rect 22972 20644 22996 20646
rect 22756 20624 23052 20644
rect 25756 20700 26052 20720
rect 25812 20698 25836 20700
rect 25892 20698 25916 20700
rect 25972 20698 25996 20700
rect 25834 20646 25836 20698
rect 25898 20646 25910 20698
rect 25972 20646 25974 20698
rect 25812 20644 25836 20646
rect 25892 20644 25916 20646
rect 25972 20644 25996 20646
rect 25756 20624 26052 20644
rect 24256 20156 24552 20176
rect 24312 20154 24336 20156
rect 24392 20154 24416 20156
rect 24472 20154 24496 20156
rect 24334 20102 24336 20154
rect 24398 20102 24410 20154
rect 24472 20102 24474 20154
rect 24312 20100 24336 20102
rect 24392 20100 24416 20102
rect 24472 20100 24496 20102
rect 24256 20080 24552 20100
rect 27256 20156 27552 20176
rect 27312 20154 27336 20156
rect 27392 20154 27416 20156
rect 27472 20154 27496 20156
rect 27334 20102 27336 20154
rect 27398 20102 27410 20154
rect 27472 20102 27474 20154
rect 27312 20100 27336 20102
rect 27392 20100 27416 20102
rect 27472 20100 27496 20102
rect 27256 20080 27552 20100
rect 22756 19612 23052 19632
rect 22812 19610 22836 19612
rect 22892 19610 22916 19612
rect 22972 19610 22996 19612
rect 22834 19558 22836 19610
rect 22898 19558 22910 19610
rect 22972 19558 22974 19610
rect 22812 19556 22836 19558
rect 22892 19556 22916 19558
rect 22972 19556 22996 19558
rect 22756 19536 23052 19556
rect 25756 19612 26052 19632
rect 25812 19610 25836 19612
rect 25892 19610 25916 19612
rect 25972 19610 25996 19612
rect 25834 19558 25836 19610
rect 25898 19558 25910 19610
rect 25972 19558 25974 19610
rect 25812 19556 25836 19558
rect 25892 19556 25916 19558
rect 25972 19556 25996 19558
rect 25756 19536 26052 19556
rect 24256 19068 24552 19088
rect 24312 19066 24336 19068
rect 24392 19066 24416 19068
rect 24472 19066 24496 19068
rect 24334 19014 24336 19066
rect 24398 19014 24410 19066
rect 24472 19014 24474 19066
rect 24312 19012 24336 19014
rect 24392 19012 24416 19014
rect 24472 19012 24496 19014
rect 24256 18992 24552 19012
rect 27256 19068 27552 19088
rect 27312 19066 27336 19068
rect 27392 19066 27416 19068
rect 27472 19066 27496 19068
rect 27334 19014 27336 19066
rect 27398 19014 27410 19066
rect 27472 19014 27474 19066
rect 27312 19012 27336 19014
rect 27392 19012 27416 19014
rect 27472 19012 27496 19014
rect 27256 18992 27552 19012
rect 22756 18524 23052 18544
rect 22812 18522 22836 18524
rect 22892 18522 22916 18524
rect 22972 18522 22996 18524
rect 22834 18470 22836 18522
rect 22898 18470 22910 18522
rect 22972 18470 22974 18522
rect 22812 18468 22836 18470
rect 22892 18468 22916 18470
rect 22972 18468 22996 18470
rect 22756 18448 23052 18468
rect 25756 18524 26052 18544
rect 25812 18522 25836 18524
rect 25892 18522 25916 18524
rect 25972 18522 25996 18524
rect 25834 18470 25836 18522
rect 25898 18470 25910 18522
rect 25972 18470 25974 18522
rect 25812 18468 25836 18470
rect 25892 18468 25916 18470
rect 25972 18468 25996 18470
rect 25756 18448 26052 18468
rect 24256 17980 24552 18000
rect 24312 17978 24336 17980
rect 24392 17978 24416 17980
rect 24472 17978 24496 17980
rect 24334 17926 24336 17978
rect 24398 17926 24410 17978
rect 24472 17926 24474 17978
rect 24312 17924 24336 17926
rect 24392 17924 24416 17926
rect 24472 17924 24496 17926
rect 24256 17904 24552 17924
rect 27256 17980 27552 18000
rect 27312 17978 27336 17980
rect 27392 17978 27416 17980
rect 27472 17978 27496 17980
rect 27334 17926 27336 17978
rect 27398 17926 27410 17978
rect 27472 17926 27474 17978
rect 27312 17924 27336 17926
rect 27392 17924 27416 17926
rect 27472 17924 27496 17926
rect 27256 17904 27552 17924
rect 22756 17436 23052 17456
rect 22812 17434 22836 17436
rect 22892 17434 22916 17436
rect 22972 17434 22996 17436
rect 22834 17382 22836 17434
rect 22898 17382 22910 17434
rect 22972 17382 22974 17434
rect 22812 17380 22836 17382
rect 22892 17380 22916 17382
rect 22972 17380 22996 17382
rect 22756 17360 23052 17380
rect 25756 17436 26052 17456
rect 25812 17434 25836 17436
rect 25892 17434 25916 17436
rect 25972 17434 25996 17436
rect 25834 17382 25836 17434
rect 25898 17382 25910 17434
rect 25972 17382 25974 17434
rect 25812 17380 25836 17382
rect 25892 17380 25916 17382
rect 25972 17380 25996 17382
rect 25756 17360 26052 17380
rect 24256 16892 24552 16912
rect 24312 16890 24336 16892
rect 24392 16890 24416 16892
rect 24472 16890 24496 16892
rect 24334 16838 24336 16890
rect 24398 16838 24410 16890
rect 24472 16838 24474 16890
rect 24312 16836 24336 16838
rect 24392 16836 24416 16838
rect 24472 16836 24496 16838
rect 24256 16816 24552 16836
rect 27256 16892 27552 16912
rect 27312 16890 27336 16892
rect 27392 16890 27416 16892
rect 27472 16890 27496 16892
rect 27334 16838 27336 16890
rect 27398 16838 27410 16890
rect 27472 16838 27474 16890
rect 27312 16836 27336 16838
rect 27392 16836 27416 16838
rect 27472 16836 27496 16838
rect 27256 16816 27552 16836
rect 22756 16348 23052 16368
rect 22812 16346 22836 16348
rect 22892 16346 22916 16348
rect 22972 16346 22996 16348
rect 22834 16294 22836 16346
rect 22898 16294 22910 16346
rect 22972 16294 22974 16346
rect 22812 16292 22836 16294
rect 22892 16292 22916 16294
rect 22972 16292 22996 16294
rect 22756 16272 23052 16292
rect 25756 16348 26052 16368
rect 25812 16346 25836 16348
rect 25892 16346 25916 16348
rect 25972 16346 25996 16348
rect 25834 16294 25836 16346
rect 25898 16294 25910 16346
rect 25972 16294 25974 16346
rect 25812 16292 25836 16294
rect 25892 16292 25916 16294
rect 25972 16292 25996 16294
rect 25756 16272 26052 16292
rect 24256 15804 24552 15824
rect 24312 15802 24336 15804
rect 24392 15802 24416 15804
rect 24472 15802 24496 15804
rect 24334 15750 24336 15802
rect 24398 15750 24410 15802
rect 24472 15750 24474 15802
rect 24312 15748 24336 15750
rect 24392 15748 24416 15750
rect 24472 15748 24496 15750
rect 24256 15728 24552 15748
rect 27256 15804 27552 15824
rect 27312 15802 27336 15804
rect 27392 15802 27416 15804
rect 27472 15802 27496 15804
rect 27334 15750 27336 15802
rect 27398 15750 27410 15802
rect 27472 15750 27474 15802
rect 27312 15748 27336 15750
rect 27392 15748 27416 15750
rect 27472 15748 27496 15750
rect 27256 15728 27552 15748
rect 22756 15260 23052 15280
rect 22812 15258 22836 15260
rect 22892 15258 22916 15260
rect 22972 15258 22996 15260
rect 22834 15206 22836 15258
rect 22898 15206 22910 15258
rect 22972 15206 22974 15258
rect 22812 15204 22836 15206
rect 22892 15204 22916 15206
rect 22972 15204 22996 15206
rect 22756 15184 23052 15204
rect 25756 15260 26052 15280
rect 25812 15258 25836 15260
rect 25892 15258 25916 15260
rect 25972 15258 25996 15260
rect 25834 15206 25836 15258
rect 25898 15206 25910 15258
rect 25972 15206 25974 15258
rect 25812 15204 25836 15206
rect 25892 15204 25916 15206
rect 25972 15204 25996 15206
rect 25756 15184 26052 15204
rect 24256 14716 24552 14736
rect 24312 14714 24336 14716
rect 24392 14714 24416 14716
rect 24472 14714 24496 14716
rect 24334 14662 24336 14714
rect 24398 14662 24410 14714
rect 24472 14662 24474 14714
rect 24312 14660 24336 14662
rect 24392 14660 24416 14662
rect 24472 14660 24496 14662
rect 24256 14640 24552 14660
rect 27256 14716 27552 14736
rect 27312 14714 27336 14716
rect 27392 14714 27416 14716
rect 27472 14714 27496 14716
rect 27334 14662 27336 14714
rect 27398 14662 27410 14714
rect 27472 14662 27474 14714
rect 27312 14660 27336 14662
rect 27392 14660 27416 14662
rect 27472 14660 27496 14662
rect 27256 14640 27552 14660
rect 22756 14172 23052 14192
rect 22812 14170 22836 14172
rect 22892 14170 22916 14172
rect 22972 14170 22996 14172
rect 22834 14118 22836 14170
rect 22898 14118 22910 14170
rect 22972 14118 22974 14170
rect 22812 14116 22836 14118
rect 22892 14116 22916 14118
rect 22972 14116 22996 14118
rect 22756 14096 23052 14116
rect 25756 14172 26052 14192
rect 25812 14170 25836 14172
rect 25892 14170 25916 14172
rect 25972 14170 25996 14172
rect 25834 14118 25836 14170
rect 25898 14118 25910 14170
rect 25972 14118 25974 14170
rect 25812 14116 25836 14118
rect 25892 14116 25916 14118
rect 25972 14116 25996 14118
rect 25756 14096 26052 14116
rect 21652 13786 21772 13814
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21256 13628 21552 13648
rect 21312 13626 21336 13628
rect 21392 13626 21416 13628
rect 21472 13626 21496 13628
rect 21334 13574 21336 13626
rect 21398 13574 21410 13626
rect 21472 13574 21474 13626
rect 21312 13572 21336 13574
rect 21392 13572 21416 13574
rect 21472 13572 21496 13574
rect 21256 13552 21552 13572
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20916 12986 20944 13398
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19338 11792 19394 11801
rect 19248 11756 19300 11762
rect 19432 11756 19484 11762
rect 19394 11736 19432 11744
rect 19338 11727 19432 11736
rect 19352 11716 19432 11727
rect 19248 11698 19300 11704
rect 19432 11698 19484 11704
rect 19260 11354 19288 11698
rect 19536 11506 19564 12174
rect 19756 11996 20052 12016
rect 19812 11994 19836 11996
rect 19892 11994 19916 11996
rect 19972 11994 19996 11996
rect 19834 11942 19836 11994
rect 19898 11942 19910 11994
rect 19972 11942 19974 11994
rect 19812 11940 19836 11942
rect 19892 11940 19916 11942
rect 19972 11940 19996 11942
rect 19756 11920 20052 11940
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19444 11478 19564 11506
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19076 9586 19104 9862
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18892 8498 18920 8978
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18984 7206 19012 9454
rect 19076 8090 19104 9522
rect 19168 8974 19196 10950
rect 19260 10742 19288 11290
rect 19444 10810 19472 11478
rect 19812 11354 19840 11562
rect 20352 11552 20404 11558
rect 20352 11494 20404 11500
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19536 10266 19564 11290
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19628 10810 19656 11154
rect 20364 11014 20392 11494
rect 20916 11150 20944 11630
rect 21008 11626 21036 12582
rect 21256 12540 21552 12560
rect 21312 12538 21336 12540
rect 21392 12538 21416 12540
rect 21472 12538 21496 12540
rect 21334 12486 21336 12538
rect 21398 12486 21410 12538
rect 21472 12486 21474 12538
rect 21312 12484 21336 12486
rect 21392 12484 21416 12486
rect 21472 12484 21496 12486
rect 21256 12464 21552 12484
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20352 11008 20404 11014
rect 20352 10950 20404 10956
rect 19756 10908 20052 10928
rect 19812 10906 19836 10908
rect 19892 10906 19916 10908
rect 19972 10906 19996 10908
rect 19834 10854 19836 10906
rect 19898 10854 19910 10906
rect 19972 10854 19974 10906
rect 19812 10852 19836 10854
rect 19892 10852 19916 10854
rect 19972 10852 19996 10854
rect 19756 10832 20052 10852
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 20088 10130 20116 10542
rect 20916 10198 20944 10610
rect 21008 10606 21036 11562
rect 21100 11354 21128 12038
rect 21256 11452 21552 11472
rect 21312 11450 21336 11452
rect 21392 11450 21416 11452
rect 21472 11450 21496 11452
rect 21334 11398 21336 11450
rect 21398 11398 21410 11450
rect 21472 11398 21474 11450
rect 21312 11396 21336 11398
rect 21392 11396 21416 11398
rect 21472 11396 21496 11398
rect 21256 11376 21552 11396
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21192 10266 21220 11018
rect 21652 10554 21680 13670
rect 21744 12986 21772 13786
rect 24256 13628 24552 13648
rect 24312 13626 24336 13628
rect 24392 13626 24416 13628
rect 24472 13626 24496 13628
rect 24334 13574 24336 13626
rect 24398 13574 24410 13626
rect 24472 13574 24474 13626
rect 24312 13572 24336 13574
rect 24392 13572 24416 13574
rect 24472 13572 24496 13574
rect 24256 13552 24552 13572
rect 27256 13628 27552 13648
rect 27312 13626 27336 13628
rect 27392 13626 27416 13628
rect 27472 13626 27496 13628
rect 27334 13574 27336 13626
rect 27398 13574 27410 13626
rect 27472 13574 27474 13626
rect 27312 13572 27336 13574
rect 27392 13572 27416 13574
rect 27472 13572 27496 13574
rect 27256 13552 27552 13572
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 22296 12918 22324 13262
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12306 22232 12786
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21744 11762 21772 12174
rect 22296 11880 22324 12854
rect 22480 12850 22508 13126
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22572 12714 22600 13194
rect 22756 13084 23052 13104
rect 22812 13082 22836 13084
rect 22892 13082 22916 13084
rect 22972 13082 22996 13084
rect 22834 13030 22836 13082
rect 22898 13030 22910 13082
rect 22972 13030 22974 13082
rect 22812 13028 22836 13030
rect 22892 13028 22916 13030
rect 22972 13028 22996 13030
rect 22756 13008 23052 13028
rect 23124 12986 23152 13194
rect 23952 12986 23980 13194
rect 25756 13084 26052 13104
rect 25812 13082 25836 13084
rect 25892 13082 25916 13084
rect 25972 13082 25996 13084
rect 25834 13030 25836 13082
rect 25898 13030 25910 13082
rect 25972 13030 25974 13082
rect 25812 13028 25836 13030
rect 25892 13028 25916 13030
rect 25972 13028 25996 13030
rect 25756 13008 26052 13028
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22572 12442 22600 12650
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22560 12164 22612 12170
rect 22664 12152 22692 12718
rect 23952 12306 23980 12922
rect 24256 12540 24552 12560
rect 24312 12538 24336 12540
rect 24392 12538 24416 12540
rect 24472 12538 24496 12540
rect 24334 12486 24336 12538
rect 24398 12486 24410 12538
rect 24472 12486 24474 12538
rect 24312 12484 24336 12486
rect 24392 12484 24416 12486
rect 24472 12484 24496 12486
rect 24256 12464 24552 12484
rect 27256 12540 27552 12560
rect 27312 12538 27336 12540
rect 27392 12538 27416 12540
rect 27472 12538 27496 12540
rect 27334 12486 27336 12538
rect 27398 12486 27410 12538
rect 27472 12486 27474 12538
rect 27312 12484 27336 12486
rect 27392 12484 27416 12486
rect 27472 12484 27496 12486
rect 27256 12464 27552 12484
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 22612 12124 22692 12152
rect 23478 12200 23534 12209
rect 23478 12135 23534 12144
rect 22560 12106 22612 12112
rect 22572 11898 22600 12106
rect 23492 12102 23520 12135
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 22756 11996 23052 12016
rect 22812 11994 22836 11996
rect 22892 11994 22916 11996
rect 22972 11994 22996 11996
rect 22834 11942 22836 11994
rect 22898 11942 22910 11994
rect 22972 11942 22974 11994
rect 24320 11966 24348 12038
rect 25756 11996 26052 12016
rect 25812 11994 25836 11996
rect 25892 11994 25916 11996
rect 25972 11994 25996 11996
rect 22812 11940 22836 11942
rect 22892 11940 22916 11942
rect 22972 11940 22996 11942
rect 22756 11920 23052 11940
rect 24308 11960 24360 11966
rect 25834 11942 25836 11994
rect 25898 11942 25910 11994
rect 25972 11942 25974 11994
rect 25812 11940 25836 11942
rect 25892 11940 25916 11942
rect 25972 11940 25996 11942
rect 25756 11920 26052 11940
rect 24308 11902 24360 11908
rect 22112 11852 22324 11880
rect 22560 11892 22612 11898
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21836 11218 21864 11630
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21744 10674 21772 11086
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21916 10600 21968 10606
rect 21652 10526 21864 10554
rect 21916 10542 21968 10548
rect 22112 10554 22140 11852
rect 22560 11834 22612 11840
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22296 11558 22324 11698
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22296 11218 22324 11494
rect 24256 11452 24552 11472
rect 24312 11450 24336 11452
rect 24392 11450 24416 11452
rect 24472 11450 24496 11452
rect 24334 11398 24336 11450
rect 24398 11398 24410 11450
rect 24472 11398 24474 11450
rect 24312 11396 24336 11398
rect 24392 11396 24416 11398
rect 24472 11396 24496 11398
rect 24256 11376 24552 11396
rect 27256 11452 27552 11472
rect 27312 11450 27336 11452
rect 27392 11450 27416 11452
rect 27472 11450 27496 11452
rect 27334 11398 27336 11450
rect 27398 11398 27410 11450
rect 27472 11398 27474 11450
rect 27312 11396 27336 11398
rect 27392 11396 27416 11398
rect 27472 11396 27496 11398
rect 27256 11376 27552 11396
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22296 10810 22324 11154
rect 28736 11121 28764 11630
rect 28722 11112 28778 11121
rect 22468 11076 22520 11082
rect 28722 11047 28778 11056
rect 22468 11018 22520 11024
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21256 10364 21552 10384
rect 21312 10362 21336 10364
rect 21392 10362 21416 10364
rect 21472 10362 21496 10364
rect 21334 10310 21336 10362
rect 21398 10310 21410 10362
rect 21472 10310 21474 10362
rect 21312 10308 21336 10310
rect 21392 10308 21416 10310
rect 21472 10308 21496 10310
rect 21256 10288 21552 10308
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 20536 10192 20588 10198
rect 20536 10134 20588 10140
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19536 9586 19564 9998
rect 20088 9926 20116 10066
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19756 9820 20052 9840
rect 19812 9818 19836 9820
rect 19892 9818 19916 9820
rect 19972 9818 19996 9820
rect 19834 9766 19836 9818
rect 19898 9766 19910 9818
rect 19972 9766 19974 9818
rect 19812 9764 19836 9766
rect 19892 9764 19916 9766
rect 19972 9764 19996 9766
rect 19756 9744 20052 9764
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19260 9178 19288 9522
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 19168 8634 19196 8910
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19168 7954 19196 8570
rect 19352 8362 19380 8842
rect 19536 8498 19564 9522
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19996 8974 20024 9386
rect 20088 9382 20116 9862
rect 20548 9450 20576 10134
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 20088 8838 20116 9318
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19756 8732 20052 8752
rect 19812 8730 19836 8732
rect 19892 8730 19916 8732
rect 19972 8730 19996 8732
rect 19834 8678 19836 8730
rect 19898 8678 19910 8730
rect 19972 8678 19974 8730
rect 19812 8676 19836 8678
rect 19892 8676 19916 8678
rect 19972 8676 19996 8678
rect 19756 8656 20052 8676
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19260 7750 19288 8230
rect 19536 7886 19564 8434
rect 19720 8022 19748 8434
rect 20088 8362 20116 8774
rect 20548 8634 20576 9386
rect 20732 8906 20760 10066
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 21100 9450 21128 9590
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21100 9042 21128 9386
rect 21256 9276 21552 9296
rect 21312 9274 21336 9276
rect 21392 9274 21416 9276
rect 21472 9274 21496 9276
rect 21334 9222 21336 9274
rect 21398 9222 21410 9274
rect 21472 9222 21474 9274
rect 21312 9220 21336 9222
rect 21392 9220 21416 9222
rect 21472 9220 21496 9222
rect 21256 9200 21552 9220
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 21652 8974 21680 10406
rect 21836 9586 21864 10526
rect 21928 9586 21956 10542
rect 22112 10526 22324 10554
rect 22112 10130 22140 10526
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22020 9722 22048 9862
rect 22112 9722 22140 9930
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21836 9330 21864 9522
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19708 8016 19760 8022
rect 19708 7958 19760 7964
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 20088 7750 20116 8298
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19260 7274 19288 7686
rect 19756 7644 20052 7664
rect 19812 7642 19836 7644
rect 19892 7642 19916 7644
rect 19972 7642 19996 7644
rect 19834 7590 19836 7642
rect 19898 7590 19910 7642
rect 19972 7590 19974 7642
rect 19812 7588 19836 7590
rect 19892 7588 19916 7590
rect 19972 7588 19996 7590
rect 19756 7568 20052 7588
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 19352 6662 19380 7278
rect 19444 6798 19472 7346
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18800 5778 18828 6122
rect 18788 5772 18840 5778
rect 18788 5714 18840 5720
rect 18892 5710 18920 6326
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18616 5370 18644 5646
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18984 5302 19012 6054
rect 19536 5914 19564 6258
rect 19628 6254 19656 7142
rect 20088 6866 20116 7686
rect 20456 7546 20484 8502
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 19756 6556 20052 6576
rect 19812 6554 19836 6556
rect 19892 6554 19916 6556
rect 19972 6554 19996 6556
rect 19834 6502 19836 6554
rect 19898 6502 19910 6554
rect 19972 6502 19974 6554
rect 19812 6500 19836 6502
rect 19892 6500 19916 6502
rect 19972 6500 19996 6502
rect 19756 6480 20052 6500
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 20076 6180 20128 6186
rect 20180 6168 20208 6598
rect 20640 6322 20668 8366
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20732 6254 20760 8842
rect 21284 8634 21312 8910
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20824 7546 20852 7958
rect 21192 7818 21220 8570
rect 21652 8498 21680 8910
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21256 8188 21552 8208
rect 21312 8186 21336 8188
rect 21392 8186 21416 8188
rect 21472 8186 21496 8188
rect 21334 8134 21336 8186
rect 21398 8134 21410 8186
rect 21472 8134 21474 8186
rect 21312 8132 21336 8134
rect 21392 8132 21416 8134
rect 21472 8132 21496 8134
rect 21256 8112 21552 8132
rect 21744 7886 21772 9318
rect 21836 9302 21956 9330
rect 21928 9110 21956 9302
rect 22112 9178 22140 9658
rect 22204 9450 22232 10406
rect 22296 9518 22324 10526
rect 22480 10470 22508 11018
rect 22756 10908 23052 10928
rect 22812 10906 22836 10908
rect 22892 10906 22916 10908
rect 22972 10906 22996 10908
rect 22834 10854 22836 10906
rect 22898 10854 22910 10906
rect 22972 10854 22974 10906
rect 22812 10852 22836 10854
rect 22892 10852 22916 10854
rect 22972 10852 22996 10854
rect 22756 10832 23052 10852
rect 25756 10908 26052 10928
rect 25812 10906 25836 10908
rect 25892 10906 25916 10908
rect 25972 10906 25996 10908
rect 25834 10854 25836 10906
rect 25898 10854 25910 10906
rect 25972 10854 25974 10906
rect 25812 10852 25836 10854
rect 25892 10852 25916 10854
rect 25972 10852 25996 10854
rect 25756 10832 26052 10852
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 21192 7478 21220 7754
rect 21744 7546 21772 7822
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21192 7002 21220 7414
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21256 7100 21552 7120
rect 21312 7098 21336 7100
rect 21392 7098 21416 7100
rect 21472 7098 21496 7100
rect 21334 7046 21336 7098
rect 21398 7046 21410 7098
rect 21472 7046 21474 7098
rect 21312 7044 21336 7046
rect 21392 7044 21416 7046
rect 21472 7044 21496 7046
rect 21256 7024 21552 7044
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 20128 6140 20208 6168
rect 20076 6122 20128 6128
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19756 5468 20052 5488
rect 19812 5466 19836 5468
rect 19892 5466 19916 5468
rect 19972 5466 19996 5468
rect 19834 5414 19836 5466
rect 19898 5414 19910 5466
rect 19972 5414 19974 5466
rect 19812 5412 19836 5414
rect 19892 5412 19916 5414
rect 19972 5412 19996 5414
rect 19756 5392 20052 5412
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18256 4924 18552 4944
rect 18312 4922 18336 4924
rect 18392 4922 18416 4924
rect 18472 4922 18496 4924
rect 18334 4870 18336 4922
rect 18398 4870 18410 4922
rect 18472 4870 18474 4922
rect 18312 4868 18336 4870
rect 18392 4868 18416 4870
rect 18472 4868 18496 4870
rect 18256 4848 18552 4868
rect 18616 4758 18644 5034
rect 18984 4826 19012 5238
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19076 4758 19104 5102
rect 19720 4826 19748 5238
rect 20180 5166 20208 6140
rect 20732 5914 20760 6190
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 20180 4826 20208 5102
rect 19708 4820 19760 4826
rect 19628 4780 19708 4808
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 18144 4684 18196 4690
rect 18144 4626 18196 4632
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18616 4214 18644 4558
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17972 3738 18000 4082
rect 18256 3836 18552 3856
rect 18312 3834 18336 3836
rect 18392 3834 18416 3836
rect 18472 3834 18496 3836
rect 18334 3782 18336 3834
rect 18398 3782 18410 3834
rect 18472 3782 18474 3834
rect 18312 3780 18336 3782
rect 18392 3780 18416 3782
rect 18472 3780 18496 3782
rect 18256 3760 18552 3780
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 16756 3292 17052 3312
rect 16812 3290 16836 3292
rect 16892 3290 16916 3292
rect 16972 3290 16996 3292
rect 16834 3238 16836 3290
rect 16898 3238 16910 3290
rect 16972 3238 16974 3290
rect 16812 3236 16836 3238
rect 16892 3236 16916 3238
rect 16972 3236 16996 3238
rect 16756 3216 17052 3236
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16960 2378 16988 2994
rect 17144 2854 17172 3402
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 3058 18000 3334
rect 18616 3194 18644 4150
rect 18892 4146 18920 4626
rect 19076 4486 19104 4694
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 19628 4282 19656 4780
rect 19708 4762 19760 4768
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20732 4758 20760 5850
rect 21008 5778 21036 6190
rect 21192 5846 21220 6734
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 6390 21680 6598
rect 21640 6384 21692 6390
rect 21640 6326 21692 6332
rect 21256 6012 21552 6032
rect 21312 6010 21336 6012
rect 21392 6010 21416 6012
rect 21472 6010 21496 6012
rect 21334 5958 21336 6010
rect 21398 5958 21410 6010
rect 21472 5958 21474 6010
rect 21312 5956 21336 5958
rect 21392 5956 21416 5958
rect 21472 5956 21496 5958
rect 21256 5936 21552 5956
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21376 5302 21404 5578
rect 21652 5370 21680 6326
rect 21744 5710 21772 7278
rect 21836 5778 21864 8570
rect 21928 6798 21956 9046
rect 22204 8906 22232 9386
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22204 8634 22232 8842
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22008 8560 22060 8566
rect 22008 8502 22060 8508
rect 22020 7954 22048 8502
rect 22296 8294 22324 8910
rect 22480 8362 22508 10406
rect 23860 10130 23888 10474
rect 24256 10364 24552 10384
rect 24312 10362 24336 10364
rect 24392 10362 24416 10364
rect 24472 10362 24496 10364
rect 24334 10310 24336 10362
rect 24398 10310 24410 10362
rect 24472 10310 24474 10362
rect 24312 10308 24336 10310
rect 24392 10308 24416 10310
rect 24472 10308 24496 10310
rect 24256 10288 24552 10308
rect 27256 10364 27552 10384
rect 27312 10362 27336 10364
rect 27392 10362 27416 10364
rect 27472 10362 27496 10364
rect 27334 10310 27336 10362
rect 27398 10310 27410 10362
rect 27472 10310 27474 10362
rect 27312 10308 27336 10310
rect 27392 10308 27416 10310
rect 27472 10308 27496 10310
rect 27256 10288 27552 10308
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 22756 9820 23052 9840
rect 22812 9818 22836 9820
rect 22892 9818 22916 9820
rect 22972 9818 22996 9820
rect 22834 9766 22836 9818
rect 22898 9766 22910 9818
rect 22972 9766 22974 9818
rect 22812 9764 22836 9766
rect 22892 9764 22916 9766
rect 22972 9764 22996 9766
rect 22756 9744 23052 9764
rect 25756 9820 26052 9840
rect 25812 9818 25836 9820
rect 25892 9818 25916 9820
rect 25972 9818 25996 9820
rect 25834 9766 25836 9818
rect 25898 9766 25910 9818
rect 25972 9766 25974 9818
rect 25812 9764 25836 9766
rect 25892 9764 25916 9766
rect 25972 9764 25996 9766
rect 25756 9744 26052 9764
rect 24256 9276 24552 9296
rect 24312 9274 24336 9276
rect 24392 9274 24416 9276
rect 24472 9274 24496 9276
rect 24334 9222 24336 9274
rect 24398 9222 24410 9274
rect 24472 9222 24474 9274
rect 24312 9220 24336 9222
rect 24392 9220 24416 9222
rect 24472 9220 24496 9222
rect 24256 9200 24552 9220
rect 27256 9276 27552 9296
rect 27312 9274 27336 9276
rect 27392 9274 27416 9276
rect 27472 9274 27496 9276
rect 27334 9222 27336 9274
rect 27398 9222 27410 9274
rect 27472 9222 27474 9274
rect 27312 9220 27336 9222
rect 27392 9220 27416 9222
rect 27472 9220 27496 9222
rect 27256 9200 27552 9220
rect 22756 8732 23052 8752
rect 22812 8730 22836 8732
rect 22892 8730 22916 8732
rect 22972 8730 22996 8732
rect 22834 8678 22836 8730
rect 22898 8678 22910 8730
rect 22972 8678 22974 8730
rect 22812 8676 22836 8678
rect 22892 8676 22916 8678
rect 22972 8676 22996 8678
rect 22756 8656 23052 8676
rect 25756 8732 26052 8752
rect 25812 8730 25836 8732
rect 25892 8730 25916 8732
rect 25972 8730 25996 8732
rect 25834 8678 25836 8730
rect 25898 8678 25910 8730
rect 25972 8678 25974 8730
rect 25812 8676 25836 8678
rect 25892 8676 25916 8678
rect 25972 8676 25996 8678
rect 25756 8656 26052 8676
rect 22468 8356 22520 8362
rect 22468 8298 22520 8304
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22296 8090 22324 8230
rect 24256 8188 24552 8208
rect 24312 8186 24336 8188
rect 24392 8186 24416 8188
rect 24472 8186 24496 8188
rect 24334 8134 24336 8186
rect 24398 8134 24410 8186
rect 24472 8134 24474 8186
rect 24312 8132 24336 8134
rect 24392 8132 24416 8134
rect 24472 8132 24496 8134
rect 24256 8112 24552 8132
rect 27256 8188 27552 8208
rect 27312 8186 27336 8188
rect 27392 8186 27416 8188
rect 27472 8186 27496 8188
rect 27334 8134 27336 8186
rect 27398 8134 27410 8186
rect 27472 8134 27474 8186
rect 27312 8132 27336 8134
rect 27392 8132 27416 8134
rect 27472 8132 27496 8134
rect 27256 8112 27552 8132
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 22756 7644 23052 7664
rect 22812 7642 22836 7644
rect 22892 7642 22916 7644
rect 22972 7642 22996 7644
rect 22834 7590 22836 7642
rect 22898 7590 22910 7642
rect 22972 7590 22974 7642
rect 22812 7588 22836 7590
rect 22892 7588 22916 7590
rect 22972 7588 22996 7590
rect 22756 7568 23052 7588
rect 25756 7644 26052 7664
rect 25812 7642 25836 7644
rect 25892 7642 25916 7644
rect 25972 7642 25996 7644
rect 25834 7590 25836 7642
rect 25898 7590 25910 7642
rect 25972 7590 25974 7642
rect 25812 7588 25836 7590
rect 25892 7588 25916 7590
rect 25972 7588 25996 7590
rect 25756 7568 26052 7588
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22020 6662 22048 7346
rect 24256 7100 24552 7120
rect 24312 7098 24336 7100
rect 24392 7098 24416 7100
rect 24472 7098 24496 7100
rect 24334 7046 24336 7098
rect 24398 7046 24410 7098
rect 24472 7046 24474 7098
rect 24312 7044 24336 7046
rect 24392 7044 24416 7046
rect 24472 7044 24496 7046
rect 24256 7024 24552 7044
rect 27256 7100 27552 7120
rect 27312 7098 27336 7100
rect 27392 7098 27416 7100
rect 27472 7098 27496 7100
rect 27334 7046 27336 7098
rect 27398 7046 27410 7098
rect 27472 7046 27474 7098
rect 27312 7044 27336 7046
rect 27392 7044 27416 7046
rect 27472 7044 27496 7046
rect 27256 7024 27552 7044
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 22020 6254 22048 6598
rect 22756 6556 23052 6576
rect 22812 6554 22836 6556
rect 22892 6554 22916 6556
rect 22972 6554 22996 6556
rect 22834 6502 22836 6554
rect 22898 6502 22910 6554
rect 22972 6502 22974 6554
rect 22812 6500 22836 6502
rect 22892 6500 22916 6502
rect 22972 6500 22996 6502
rect 22756 6480 23052 6500
rect 25756 6556 26052 6576
rect 25812 6554 25836 6556
rect 25892 6554 25916 6556
rect 25972 6554 25996 6556
rect 25834 6502 25836 6554
rect 25898 6502 25910 6554
rect 25972 6502 25974 6554
rect 25812 6500 25836 6502
rect 25892 6500 25916 6502
rect 25972 6500 25996 6502
rect 25756 6480 26052 6500
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22020 5778 22048 6190
rect 24256 6012 24552 6032
rect 24312 6010 24336 6012
rect 24392 6010 24416 6012
rect 24472 6010 24496 6012
rect 24334 5958 24336 6010
rect 24398 5958 24410 6010
rect 24472 5958 24474 6010
rect 24312 5956 24336 5958
rect 24392 5956 24416 5958
rect 24472 5956 24496 5958
rect 24256 5936 24552 5956
rect 27256 6012 27552 6032
rect 27312 6010 27336 6012
rect 27392 6010 27416 6012
rect 27472 6010 27496 6012
rect 27334 5958 27336 6010
rect 27398 5958 27410 6010
rect 27472 5958 27474 6010
rect 27312 5956 27336 5958
rect 27392 5956 27416 5958
rect 27472 5956 27496 5958
rect 27256 5936 27552 5956
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21640 5364 21692 5370
rect 21640 5306 21692 5312
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21256 4924 21552 4944
rect 21312 4922 21336 4924
rect 21392 4922 21416 4924
rect 21472 4922 21496 4924
rect 21334 4870 21336 4922
rect 21398 4870 21410 4922
rect 21472 4870 21474 4922
rect 21312 4868 21336 4870
rect 21392 4868 21416 4870
rect 21472 4868 21496 4870
rect 21256 4848 21552 4868
rect 21744 4758 21772 5646
rect 21836 5370 21864 5714
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 22020 4826 22048 5714
rect 22756 5468 23052 5488
rect 22812 5466 22836 5468
rect 22892 5466 22916 5468
rect 22972 5466 22996 5468
rect 22834 5414 22836 5466
rect 22898 5414 22910 5466
rect 22972 5414 22974 5466
rect 22812 5412 22836 5414
rect 22892 5412 22916 5414
rect 22972 5412 22996 5414
rect 22756 5392 23052 5412
rect 25756 5468 26052 5488
rect 25812 5466 25836 5468
rect 25892 5466 25916 5468
rect 25972 5466 25996 5468
rect 25834 5414 25836 5466
rect 25898 5414 25910 5466
rect 25972 5414 25974 5466
rect 25812 5412 25836 5414
rect 25892 5412 25916 5414
rect 25972 5412 25996 5414
rect 25756 5392 26052 5412
rect 24256 4924 24552 4944
rect 24312 4922 24336 4924
rect 24392 4922 24416 4924
rect 24472 4922 24496 4924
rect 24334 4870 24336 4922
rect 24398 4870 24410 4922
rect 24472 4870 24474 4922
rect 24312 4868 24336 4870
rect 24392 4868 24416 4870
rect 24472 4868 24496 4870
rect 24256 4848 24552 4868
rect 27256 4924 27552 4944
rect 27312 4922 27336 4924
rect 27392 4922 27416 4924
rect 27472 4922 27496 4924
rect 27334 4870 27336 4922
rect 27398 4870 27410 4922
rect 27472 4870 27474 4922
rect 27312 4868 27336 4870
rect 27392 4868 27416 4870
rect 27472 4868 27496 4870
rect 27256 4848 27552 4868
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 19756 4380 20052 4400
rect 19812 4378 19836 4380
rect 19892 4378 19916 4380
rect 19972 4378 19996 4380
rect 19834 4326 19836 4378
rect 19898 4326 19910 4378
rect 19972 4326 19974 4378
rect 19812 4324 19836 4326
rect 19892 4324 19916 4326
rect 19972 4324 19996 4326
rect 19756 4304 20052 4324
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19352 3738 19380 3946
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18708 3126 18736 3470
rect 19628 3398 19656 4082
rect 20180 3738 20208 4422
rect 22756 4380 23052 4400
rect 22812 4378 22836 4380
rect 22892 4378 22916 4380
rect 22972 4378 22996 4380
rect 22834 4326 22836 4378
rect 22898 4326 22910 4378
rect 22972 4326 22974 4378
rect 22812 4324 22836 4326
rect 22892 4324 22916 4326
rect 22972 4324 22996 4326
rect 22756 4304 23052 4324
rect 25756 4380 26052 4400
rect 25812 4378 25836 4380
rect 25892 4378 25916 4380
rect 25972 4378 25996 4380
rect 25834 4326 25836 4378
rect 25898 4326 25910 4378
rect 25972 4326 25974 4378
rect 25812 4324 25836 4326
rect 25892 4324 25916 4326
rect 25972 4324 25996 4326
rect 25756 4304 26052 4324
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19756 3292 20052 3312
rect 19812 3290 19836 3292
rect 19892 3290 19916 3292
rect 19972 3290 19996 3292
rect 19834 3238 19836 3290
rect 19898 3238 19910 3290
rect 19972 3238 19974 3290
rect 19812 3236 19836 3238
rect 19892 3236 19916 3238
rect 19972 3236 19996 3238
rect 19756 3216 20052 3236
rect 20456 3194 20484 3878
rect 21256 3836 21552 3856
rect 21312 3834 21336 3836
rect 21392 3834 21416 3836
rect 21472 3834 21496 3836
rect 21334 3782 21336 3834
rect 21398 3782 21410 3834
rect 21472 3782 21474 3834
rect 21312 3780 21336 3782
rect 21392 3780 21416 3782
rect 21472 3780 21496 3782
rect 21256 3760 21552 3780
rect 24256 3836 24552 3856
rect 24312 3834 24336 3836
rect 24392 3834 24416 3836
rect 24472 3834 24496 3836
rect 24334 3782 24336 3834
rect 24398 3782 24410 3834
rect 24472 3782 24474 3834
rect 24312 3780 24336 3782
rect 24392 3780 24416 3782
rect 24472 3780 24496 3782
rect 24256 3760 24552 3780
rect 27256 3836 27552 3856
rect 27312 3834 27336 3836
rect 27392 3834 27416 3836
rect 27472 3834 27496 3836
rect 27334 3782 27336 3834
rect 27398 3782 27410 3834
rect 27472 3782 27474 3834
rect 27312 3780 27336 3782
rect 27392 3780 27416 3782
rect 27472 3780 27496 3782
rect 27256 3760 27552 3780
rect 22756 3292 23052 3312
rect 22812 3290 22836 3292
rect 22892 3290 22916 3292
rect 22972 3290 22996 3292
rect 22834 3238 22836 3290
rect 22898 3238 22910 3290
rect 22972 3238 22974 3290
rect 22812 3236 22836 3238
rect 22892 3236 22916 3238
rect 22972 3236 22996 3238
rect 22756 3216 23052 3236
rect 25756 3292 26052 3312
rect 25812 3290 25836 3292
rect 25892 3290 25916 3292
rect 25972 3290 25996 3292
rect 25834 3238 25836 3290
rect 25898 3238 25910 3290
rect 25972 3238 25974 3290
rect 25812 3236 25836 3238
rect 25892 3236 25916 3238
rect 25972 3236 25996 3238
rect 25756 3216 26052 3236
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 2650 17540 2790
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17972 2582 18000 2994
rect 18256 2748 18552 2768
rect 18312 2746 18336 2748
rect 18392 2746 18416 2748
rect 18472 2746 18496 2748
rect 18334 2694 18336 2746
rect 18398 2694 18410 2746
rect 18472 2694 18474 2746
rect 18312 2692 18336 2694
rect 18392 2692 18416 2694
rect 18472 2692 18496 2694
rect 18256 2672 18552 2692
rect 21256 2748 21552 2768
rect 21312 2746 21336 2748
rect 21392 2746 21416 2748
rect 21472 2746 21496 2748
rect 21334 2694 21336 2746
rect 21398 2694 21410 2746
rect 21472 2694 21474 2746
rect 21312 2692 21336 2694
rect 21392 2692 21416 2694
rect 21472 2692 21496 2694
rect 21256 2672 21552 2692
rect 24256 2748 24552 2768
rect 24312 2746 24336 2748
rect 24392 2746 24416 2748
rect 24472 2746 24496 2748
rect 24334 2694 24336 2746
rect 24398 2694 24410 2746
rect 24472 2694 24474 2746
rect 24312 2692 24336 2694
rect 24392 2692 24416 2694
rect 24472 2692 24496 2694
rect 24256 2672 24552 2692
rect 27256 2748 27552 2768
rect 27312 2746 27336 2748
rect 27392 2746 27416 2748
rect 27472 2746 27496 2748
rect 27334 2694 27336 2746
rect 27398 2694 27410 2746
rect 27472 2694 27474 2746
rect 27312 2692 27336 2694
rect 27392 2692 27416 2694
rect 27472 2692 27496 2694
rect 27256 2672 27552 2692
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 10756 2204 11052 2224
rect 10812 2202 10836 2204
rect 10892 2202 10916 2204
rect 10972 2202 10996 2204
rect 10834 2150 10836 2202
rect 10898 2150 10910 2202
rect 10972 2150 10974 2202
rect 10812 2148 10836 2150
rect 10892 2148 10916 2150
rect 10972 2148 10996 2150
rect 10756 2128 11052 2148
rect 13756 2204 14052 2224
rect 13812 2202 13836 2204
rect 13892 2202 13916 2204
rect 13972 2202 13996 2204
rect 13834 2150 13836 2202
rect 13898 2150 13910 2202
rect 13972 2150 13974 2202
rect 13812 2148 13836 2150
rect 13892 2148 13916 2150
rect 13972 2148 13996 2150
rect 13756 2128 14052 2148
rect 16756 2204 17052 2224
rect 16812 2202 16836 2204
rect 16892 2202 16916 2204
rect 16972 2202 16996 2204
rect 16834 2150 16836 2202
rect 16898 2150 16910 2202
rect 16972 2150 16974 2202
rect 16812 2148 16836 2150
rect 16892 2148 16916 2150
rect 16972 2148 16996 2150
rect 16756 2128 17052 2148
rect 18248 82 18276 2314
rect 19756 2204 20052 2224
rect 19812 2202 19836 2204
rect 19892 2202 19916 2204
rect 19972 2202 19996 2204
rect 19834 2150 19836 2202
rect 19898 2150 19910 2202
rect 19972 2150 19974 2202
rect 19812 2148 19836 2150
rect 19892 2148 19916 2150
rect 19972 2148 19996 2150
rect 19756 2128 20052 2148
rect 22756 2204 23052 2224
rect 22812 2202 22836 2204
rect 22892 2202 22916 2204
rect 22972 2202 22996 2204
rect 22834 2150 22836 2202
rect 22898 2150 22910 2202
rect 22972 2150 22974 2202
rect 22812 2148 22836 2150
rect 22892 2148 22916 2150
rect 22972 2148 22996 2150
rect 22756 2128 23052 2148
rect 25756 2204 26052 2224
rect 25812 2202 25836 2204
rect 25892 2202 25916 2204
rect 25972 2202 25996 2204
rect 25834 2150 25836 2202
rect 25898 2150 25910 2202
rect 25972 2150 25974 2202
rect 25812 2148 25836 2150
rect 25892 2148 25916 2150
rect 25972 2148 25996 2150
rect 25756 2128 26052 2148
rect 18510 82 18566 800
rect 9956 60 10008 66
rect 9218 0 9274 54
rect 18248 54 18566 82
rect 9956 2 10008 8
rect 18510 0 18566 54
rect 27710 0 27766 800
<< via2 >>
rect 1756 29402 1812 29404
rect 1836 29402 1892 29404
rect 1916 29402 1972 29404
rect 1996 29402 2052 29404
rect 1756 29350 1782 29402
rect 1782 29350 1812 29402
rect 1836 29350 1846 29402
rect 1846 29350 1892 29402
rect 1916 29350 1962 29402
rect 1962 29350 1972 29402
rect 1996 29350 2026 29402
rect 2026 29350 2052 29402
rect 1756 29348 1812 29350
rect 1836 29348 1892 29350
rect 1916 29348 1972 29350
rect 1996 29348 2052 29350
rect 4756 29402 4812 29404
rect 4836 29402 4892 29404
rect 4916 29402 4972 29404
rect 4996 29402 5052 29404
rect 4756 29350 4782 29402
rect 4782 29350 4812 29402
rect 4836 29350 4846 29402
rect 4846 29350 4892 29402
rect 4916 29350 4962 29402
rect 4962 29350 4972 29402
rect 4996 29350 5026 29402
rect 5026 29350 5052 29402
rect 4756 29348 4812 29350
rect 4836 29348 4892 29350
rect 4916 29348 4972 29350
rect 4996 29348 5052 29350
rect 7756 29402 7812 29404
rect 7836 29402 7892 29404
rect 7916 29402 7972 29404
rect 7996 29402 8052 29404
rect 7756 29350 7782 29402
rect 7782 29350 7812 29402
rect 7836 29350 7846 29402
rect 7846 29350 7892 29402
rect 7916 29350 7962 29402
rect 7962 29350 7972 29402
rect 7996 29350 8026 29402
rect 8026 29350 8052 29402
rect 7756 29348 7812 29350
rect 7836 29348 7892 29350
rect 7916 29348 7972 29350
rect 7996 29348 8052 29350
rect 10756 29402 10812 29404
rect 10836 29402 10892 29404
rect 10916 29402 10972 29404
rect 10996 29402 11052 29404
rect 10756 29350 10782 29402
rect 10782 29350 10812 29402
rect 10836 29350 10846 29402
rect 10846 29350 10892 29402
rect 10916 29350 10962 29402
rect 10962 29350 10972 29402
rect 10996 29350 11026 29402
rect 11026 29350 11052 29402
rect 10756 29348 10812 29350
rect 10836 29348 10892 29350
rect 10916 29348 10972 29350
rect 10996 29348 11052 29350
rect 13756 29402 13812 29404
rect 13836 29402 13892 29404
rect 13916 29402 13972 29404
rect 13996 29402 14052 29404
rect 13756 29350 13782 29402
rect 13782 29350 13812 29402
rect 13836 29350 13846 29402
rect 13846 29350 13892 29402
rect 13916 29350 13962 29402
rect 13962 29350 13972 29402
rect 13996 29350 14026 29402
rect 14026 29350 14052 29402
rect 13756 29348 13812 29350
rect 13836 29348 13892 29350
rect 13916 29348 13972 29350
rect 13996 29348 14052 29350
rect 16756 29402 16812 29404
rect 16836 29402 16892 29404
rect 16916 29402 16972 29404
rect 16996 29402 17052 29404
rect 16756 29350 16782 29402
rect 16782 29350 16812 29402
rect 16836 29350 16846 29402
rect 16846 29350 16892 29402
rect 16916 29350 16962 29402
rect 16962 29350 16972 29402
rect 16996 29350 17026 29402
rect 17026 29350 17052 29402
rect 16756 29348 16812 29350
rect 16836 29348 16892 29350
rect 16916 29348 16972 29350
rect 16996 29348 17052 29350
rect 19756 29402 19812 29404
rect 19836 29402 19892 29404
rect 19916 29402 19972 29404
rect 19996 29402 20052 29404
rect 19756 29350 19782 29402
rect 19782 29350 19812 29402
rect 19836 29350 19846 29402
rect 19846 29350 19892 29402
rect 19916 29350 19962 29402
rect 19962 29350 19972 29402
rect 19996 29350 20026 29402
rect 20026 29350 20052 29402
rect 19756 29348 19812 29350
rect 19836 29348 19892 29350
rect 19916 29348 19972 29350
rect 19996 29348 20052 29350
rect 22756 29402 22812 29404
rect 22836 29402 22892 29404
rect 22916 29402 22972 29404
rect 22996 29402 23052 29404
rect 22756 29350 22782 29402
rect 22782 29350 22812 29402
rect 22836 29350 22846 29402
rect 22846 29350 22892 29402
rect 22916 29350 22962 29402
rect 22962 29350 22972 29402
rect 22996 29350 23026 29402
rect 23026 29350 23052 29402
rect 22756 29348 22812 29350
rect 22836 29348 22892 29350
rect 22916 29348 22972 29350
rect 22996 29348 23052 29350
rect 3256 28858 3312 28860
rect 3336 28858 3392 28860
rect 3416 28858 3472 28860
rect 3496 28858 3552 28860
rect 3256 28806 3282 28858
rect 3282 28806 3312 28858
rect 3336 28806 3346 28858
rect 3346 28806 3392 28858
rect 3416 28806 3462 28858
rect 3462 28806 3472 28858
rect 3496 28806 3526 28858
rect 3526 28806 3552 28858
rect 3256 28804 3312 28806
rect 3336 28804 3392 28806
rect 3416 28804 3472 28806
rect 3496 28804 3552 28806
rect 6256 28858 6312 28860
rect 6336 28858 6392 28860
rect 6416 28858 6472 28860
rect 6496 28858 6552 28860
rect 6256 28806 6282 28858
rect 6282 28806 6312 28858
rect 6336 28806 6346 28858
rect 6346 28806 6392 28858
rect 6416 28806 6462 28858
rect 6462 28806 6472 28858
rect 6496 28806 6526 28858
rect 6526 28806 6552 28858
rect 6256 28804 6312 28806
rect 6336 28804 6392 28806
rect 6416 28804 6472 28806
rect 6496 28804 6552 28806
rect 9256 28858 9312 28860
rect 9336 28858 9392 28860
rect 9416 28858 9472 28860
rect 9496 28858 9552 28860
rect 9256 28806 9282 28858
rect 9282 28806 9312 28858
rect 9336 28806 9346 28858
rect 9346 28806 9392 28858
rect 9416 28806 9462 28858
rect 9462 28806 9472 28858
rect 9496 28806 9526 28858
rect 9526 28806 9552 28858
rect 9256 28804 9312 28806
rect 9336 28804 9392 28806
rect 9416 28804 9472 28806
rect 9496 28804 9552 28806
rect 12256 28858 12312 28860
rect 12336 28858 12392 28860
rect 12416 28858 12472 28860
rect 12496 28858 12552 28860
rect 12256 28806 12282 28858
rect 12282 28806 12312 28858
rect 12336 28806 12346 28858
rect 12346 28806 12392 28858
rect 12416 28806 12462 28858
rect 12462 28806 12472 28858
rect 12496 28806 12526 28858
rect 12526 28806 12552 28858
rect 12256 28804 12312 28806
rect 12336 28804 12392 28806
rect 12416 28804 12472 28806
rect 12496 28804 12552 28806
rect 15256 28858 15312 28860
rect 15336 28858 15392 28860
rect 15416 28858 15472 28860
rect 15496 28858 15552 28860
rect 15256 28806 15282 28858
rect 15282 28806 15312 28858
rect 15336 28806 15346 28858
rect 15346 28806 15392 28858
rect 15416 28806 15462 28858
rect 15462 28806 15472 28858
rect 15496 28806 15526 28858
rect 15526 28806 15552 28858
rect 15256 28804 15312 28806
rect 15336 28804 15392 28806
rect 15416 28804 15472 28806
rect 15496 28804 15552 28806
rect 18256 28858 18312 28860
rect 18336 28858 18392 28860
rect 18416 28858 18472 28860
rect 18496 28858 18552 28860
rect 18256 28806 18282 28858
rect 18282 28806 18312 28858
rect 18336 28806 18346 28858
rect 18346 28806 18392 28858
rect 18416 28806 18462 28858
rect 18462 28806 18472 28858
rect 18496 28806 18526 28858
rect 18526 28806 18552 28858
rect 18256 28804 18312 28806
rect 18336 28804 18392 28806
rect 18416 28804 18472 28806
rect 18496 28804 18552 28806
rect 21256 28858 21312 28860
rect 21336 28858 21392 28860
rect 21416 28858 21472 28860
rect 21496 28858 21552 28860
rect 21256 28806 21282 28858
rect 21282 28806 21312 28858
rect 21336 28806 21346 28858
rect 21346 28806 21392 28858
rect 21416 28806 21462 28858
rect 21462 28806 21472 28858
rect 21496 28806 21526 28858
rect 21526 28806 21552 28858
rect 21256 28804 21312 28806
rect 21336 28804 21392 28806
rect 21416 28804 21472 28806
rect 21496 28804 21552 28806
rect 24256 28858 24312 28860
rect 24336 28858 24392 28860
rect 24416 28858 24472 28860
rect 24496 28858 24552 28860
rect 24256 28806 24282 28858
rect 24282 28806 24312 28858
rect 24336 28806 24346 28858
rect 24346 28806 24392 28858
rect 24416 28806 24462 28858
rect 24462 28806 24472 28858
rect 24496 28806 24526 28858
rect 24526 28806 24552 28858
rect 24256 28804 24312 28806
rect 24336 28804 24392 28806
rect 24416 28804 24472 28806
rect 24496 28804 24552 28806
rect 1756 28314 1812 28316
rect 1836 28314 1892 28316
rect 1916 28314 1972 28316
rect 1996 28314 2052 28316
rect 1756 28262 1782 28314
rect 1782 28262 1812 28314
rect 1836 28262 1846 28314
rect 1846 28262 1892 28314
rect 1916 28262 1962 28314
rect 1962 28262 1972 28314
rect 1996 28262 2026 28314
rect 2026 28262 2052 28314
rect 1756 28260 1812 28262
rect 1836 28260 1892 28262
rect 1916 28260 1972 28262
rect 1996 28260 2052 28262
rect 4756 28314 4812 28316
rect 4836 28314 4892 28316
rect 4916 28314 4972 28316
rect 4996 28314 5052 28316
rect 4756 28262 4782 28314
rect 4782 28262 4812 28314
rect 4836 28262 4846 28314
rect 4846 28262 4892 28314
rect 4916 28262 4962 28314
rect 4962 28262 4972 28314
rect 4996 28262 5026 28314
rect 5026 28262 5052 28314
rect 4756 28260 4812 28262
rect 4836 28260 4892 28262
rect 4916 28260 4972 28262
rect 4996 28260 5052 28262
rect 7756 28314 7812 28316
rect 7836 28314 7892 28316
rect 7916 28314 7972 28316
rect 7996 28314 8052 28316
rect 7756 28262 7782 28314
rect 7782 28262 7812 28314
rect 7836 28262 7846 28314
rect 7846 28262 7892 28314
rect 7916 28262 7962 28314
rect 7962 28262 7972 28314
rect 7996 28262 8026 28314
rect 8026 28262 8052 28314
rect 7756 28260 7812 28262
rect 7836 28260 7892 28262
rect 7916 28260 7972 28262
rect 7996 28260 8052 28262
rect 10756 28314 10812 28316
rect 10836 28314 10892 28316
rect 10916 28314 10972 28316
rect 10996 28314 11052 28316
rect 10756 28262 10782 28314
rect 10782 28262 10812 28314
rect 10836 28262 10846 28314
rect 10846 28262 10892 28314
rect 10916 28262 10962 28314
rect 10962 28262 10972 28314
rect 10996 28262 11026 28314
rect 11026 28262 11052 28314
rect 10756 28260 10812 28262
rect 10836 28260 10892 28262
rect 10916 28260 10972 28262
rect 10996 28260 11052 28262
rect 13756 28314 13812 28316
rect 13836 28314 13892 28316
rect 13916 28314 13972 28316
rect 13996 28314 14052 28316
rect 13756 28262 13782 28314
rect 13782 28262 13812 28314
rect 13836 28262 13846 28314
rect 13846 28262 13892 28314
rect 13916 28262 13962 28314
rect 13962 28262 13972 28314
rect 13996 28262 14026 28314
rect 14026 28262 14052 28314
rect 13756 28260 13812 28262
rect 13836 28260 13892 28262
rect 13916 28260 13972 28262
rect 13996 28260 14052 28262
rect 16756 28314 16812 28316
rect 16836 28314 16892 28316
rect 16916 28314 16972 28316
rect 16996 28314 17052 28316
rect 16756 28262 16782 28314
rect 16782 28262 16812 28314
rect 16836 28262 16846 28314
rect 16846 28262 16892 28314
rect 16916 28262 16962 28314
rect 16962 28262 16972 28314
rect 16996 28262 17026 28314
rect 17026 28262 17052 28314
rect 16756 28260 16812 28262
rect 16836 28260 16892 28262
rect 16916 28260 16972 28262
rect 16996 28260 17052 28262
rect 19756 28314 19812 28316
rect 19836 28314 19892 28316
rect 19916 28314 19972 28316
rect 19996 28314 20052 28316
rect 19756 28262 19782 28314
rect 19782 28262 19812 28314
rect 19836 28262 19846 28314
rect 19846 28262 19892 28314
rect 19916 28262 19962 28314
rect 19962 28262 19972 28314
rect 19996 28262 20026 28314
rect 20026 28262 20052 28314
rect 19756 28260 19812 28262
rect 19836 28260 19892 28262
rect 19916 28260 19972 28262
rect 19996 28260 20052 28262
rect 22756 28314 22812 28316
rect 22836 28314 22892 28316
rect 22916 28314 22972 28316
rect 22996 28314 23052 28316
rect 22756 28262 22782 28314
rect 22782 28262 22812 28314
rect 22836 28262 22846 28314
rect 22846 28262 22892 28314
rect 22916 28262 22962 28314
rect 22962 28262 22972 28314
rect 22996 28262 23026 28314
rect 23026 28262 23052 28314
rect 22756 28260 22812 28262
rect 22836 28260 22892 28262
rect 22916 28260 22972 28262
rect 22996 28260 23052 28262
rect 3256 27770 3312 27772
rect 3336 27770 3392 27772
rect 3416 27770 3472 27772
rect 3496 27770 3552 27772
rect 3256 27718 3282 27770
rect 3282 27718 3312 27770
rect 3336 27718 3346 27770
rect 3346 27718 3392 27770
rect 3416 27718 3462 27770
rect 3462 27718 3472 27770
rect 3496 27718 3526 27770
rect 3526 27718 3552 27770
rect 3256 27716 3312 27718
rect 3336 27716 3392 27718
rect 3416 27716 3472 27718
rect 3496 27716 3552 27718
rect 6256 27770 6312 27772
rect 6336 27770 6392 27772
rect 6416 27770 6472 27772
rect 6496 27770 6552 27772
rect 6256 27718 6282 27770
rect 6282 27718 6312 27770
rect 6336 27718 6346 27770
rect 6346 27718 6392 27770
rect 6416 27718 6462 27770
rect 6462 27718 6472 27770
rect 6496 27718 6526 27770
rect 6526 27718 6552 27770
rect 6256 27716 6312 27718
rect 6336 27716 6392 27718
rect 6416 27716 6472 27718
rect 6496 27716 6552 27718
rect 9256 27770 9312 27772
rect 9336 27770 9392 27772
rect 9416 27770 9472 27772
rect 9496 27770 9552 27772
rect 9256 27718 9282 27770
rect 9282 27718 9312 27770
rect 9336 27718 9346 27770
rect 9346 27718 9392 27770
rect 9416 27718 9462 27770
rect 9462 27718 9472 27770
rect 9496 27718 9526 27770
rect 9526 27718 9552 27770
rect 9256 27716 9312 27718
rect 9336 27716 9392 27718
rect 9416 27716 9472 27718
rect 9496 27716 9552 27718
rect 12256 27770 12312 27772
rect 12336 27770 12392 27772
rect 12416 27770 12472 27772
rect 12496 27770 12552 27772
rect 12256 27718 12282 27770
rect 12282 27718 12312 27770
rect 12336 27718 12346 27770
rect 12346 27718 12392 27770
rect 12416 27718 12462 27770
rect 12462 27718 12472 27770
rect 12496 27718 12526 27770
rect 12526 27718 12552 27770
rect 12256 27716 12312 27718
rect 12336 27716 12392 27718
rect 12416 27716 12472 27718
rect 12496 27716 12552 27718
rect 15256 27770 15312 27772
rect 15336 27770 15392 27772
rect 15416 27770 15472 27772
rect 15496 27770 15552 27772
rect 15256 27718 15282 27770
rect 15282 27718 15312 27770
rect 15336 27718 15346 27770
rect 15346 27718 15392 27770
rect 15416 27718 15462 27770
rect 15462 27718 15472 27770
rect 15496 27718 15526 27770
rect 15526 27718 15552 27770
rect 15256 27716 15312 27718
rect 15336 27716 15392 27718
rect 15416 27716 15472 27718
rect 15496 27716 15552 27718
rect 18256 27770 18312 27772
rect 18336 27770 18392 27772
rect 18416 27770 18472 27772
rect 18496 27770 18552 27772
rect 18256 27718 18282 27770
rect 18282 27718 18312 27770
rect 18336 27718 18346 27770
rect 18346 27718 18392 27770
rect 18416 27718 18462 27770
rect 18462 27718 18472 27770
rect 18496 27718 18526 27770
rect 18526 27718 18552 27770
rect 18256 27716 18312 27718
rect 18336 27716 18392 27718
rect 18416 27716 18472 27718
rect 18496 27716 18552 27718
rect 21256 27770 21312 27772
rect 21336 27770 21392 27772
rect 21416 27770 21472 27772
rect 21496 27770 21552 27772
rect 21256 27718 21282 27770
rect 21282 27718 21312 27770
rect 21336 27718 21346 27770
rect 21346 27718 21392 27770
rect 21416 27718 21462 27770
rect 21462 27718 21472 27770
rect 21496 27718 21526 27770
rect 21526 27718 21552 27770
rect 21256 27716 21312 27718
rect 21336 27716 21392 27718
rect 21416 27716 21472 27718
rect 21496 27716 21552 27718
rect 24256 27770 24312 27772
rect 24336 27770 24392 27772
rect 24416 27770 24472 27772
rect 24496 27770 24552 27772
rect 24256 27718 24282 27770
rect 24282 27718 24312 27770
rect 24336 27718 24346 27770
rect 24346 27718 24392 27770
rect 24416 27718 24462 27770
rect 24462 27718 24472 27770
rect 24496 27718 24526 27770
rect 24526 27718 24552 27770
rect 24256 27716 24312 27718
rect 24336 27716 24392 27718
rect 24416 27716 24472 27718
rect 24496 27716 24552 27718
rect 25756 29402 25812 29404
rect 25836 29402 25892 29404
rect 25916 29402 25972 29404
rect 25996 29402 26052 29404
rect 25756 29350 25782 29402
rect 25782 29350 25812 29402
rect 25836 29350 25846 29402
rect 25846 29350 25892 29402
rect 25916 29350 25962 29402
rect 25962 29350 25972 29402
rect 25996 29350 26026 29402
rect 26026 29350 26052 29402
rect 25756 29348 25812 29350
rect 25836 29348 25892 29350
rect 25916 29348 25972 29350
rect 25996 29348 26052 29350
rect 27256 28858 27312 28860
rect 27336 28858 27392 28860
rect 27416 28858 27472 28860
rect 27496 28858 27552 28860
rect 27256 28806 27282 28858
rect 27282 28806 27312 28858
rect 27336 28806 27346 28858
rect 27346 28806 27392 28858
rect 27416 28806 27462 28858
rect 27462 28806 27472 28858
rect 27496 28806 27526 28858
rect 27526 28806 27552 28858
rect 27256 28804 27312 28806
rect 27336 28804 27392 28806
rect 27416 28804 27472 28806
rect 27496 28804 27552 28806
rect 25756 28314 25812 28316
rect 25836 28314 25892 28316
rect 25916 28314 25972 28316
rect 25996 28314 26052 28316
rect 25756 28262 25782 28314
rect 25782 28262 25812 28314
rect 25836 28262 25846 28314
rect 25846 28262 25892 28314
rect 25916 28262 25962 28314
rect 25962 28262 25972 28314
rect 25996 28262 26026 28314
rect 26026 28262 26052 28314
rect 25756 28260 25812 28262
rect 25836 28260 25892 28262
rect 25916 28260 25972 28262
rect 25996 28260 26052 28262
rect 27256 27770 27312 27772
rect 27336 27770 27392 27772
rect 27416 27770 27472 27772
rect 27496 27770 27552 27772
rect 27256 27718 27282 27770
rect 27282 27718 27312 27770
rect 27336 27718 27346 27770
rect 27346 27718 27392 27770
rect 27416 27718 27462 27770
rect 27462 27718 27472 27770
rect 27496 27718 27526 27770
rect 27526 27718 27552 27770
rect 27256 27716 27312 27718
rect 27336 27716 27392 27718
rect 27416 27716 27472 27718
rect 27496 27716 27552 27718
rect 1756 27226 1812 27228
rect 1836 27226 1892 27228
rect 1916 27226 1972 27228
rect 1996 27226 2052 27228
rect 1756 27174 1782 27226
rect 1782 27174 1812 27226
rect 1836 27174 1846 27226
rect 1846 27174 1892 27226
rect 1916 27174 1962 27226
rect 1962 27174 1972 27226
rect 1996 27174 2026 27226
rect 2026 27174 2052 27226
rect 1756 27172 1812 27174
rect 1836 27172 1892 27174
rect 1916 27172 1972 27174
rect 1996 27172 2052 27174
rect 4756 27226 4812 27228
rect 4836 27226 4892 27228
rect 4916 27226 4972 27228
rect 4996 27226 5052 27228
rect 4756 27174 4782 27226
rect 4782 27174 4812 27226
rect 4836 27174 4846 27226
rect 4846 27174 4892 27226
rect 4916 27174 4962 27226
rect 4962 27174 4972 27226
rect 4996 27174 5026 27226
rect 5026 27174 5052 27226
rect 4756 27172 4812 27174
rect 4836 27172 4892 27174
rect 4916 27172 4972 27174
rect 4996 27172 5052 27174
rect 7756 27226 7812 27228
rect 7836 27226 7892 27228
rect 7916 27226 7972 27228
rect 7996 27226 8052 27228
rect 7756 27174 7782 27226
rect 7782 27174 7812 27226
rect 7836 27174 7846 27226
rect 7846 27174 7892 27226
rect 7916 27174 7962 27226
rect 7962 27174 7972 27226
rect 7996 27174 8026 27226
rect 8026 27174 8052 27226
rect 7756 27172 7812 27174
rect 7836 27172 7892 27174
rect 7916 27172 7972 27174
rect 7996 27172 8052 27174
rect 10756 27226 10812 27228
rect 10836 27226 10892 27228
rect 10916 27226 10972 27228
rect 10996 27226 11052 27228
rect 10756 27174 10782 27226
rect 10782 27174 10812 27226
rect 10836 27174 10846 27226
rect 10846 27174 10892 27226
rect 10916 27174 10962 27226
rect 10962 27174 10972 27226
rect 10996 27174 11026 27226
rect 11026 27174 11052 27226
rect 10756 27172 10812 27174
rect 10836 27172 10892 27174
rect 10916 27172 10972 27174
rect 10996 27172 11052 27174
rect 13756 27226 13812 27228
rect 13836 27226 13892 27228
rect 13916 27226 13972 27228
rect 13996 27226 14052 27228
rect 13756 27174 13782 27226
rect 13782 27174 13812 27226
rect 13836 27174 13846 27226
rect 13846 27174 13892 27226
rect 13916 27174 13962 27226
rect 13962 27174 13972 27226
rect 13996 27174 14026 27226
rect 14026 27174 14052 27226
rect 13756 27172 13812 27174
rect 13836 27172 13892 27174
rect 13916 27172 13972 27174
rect 13996 27172 14052 27174
rect 16756 27226 16812 27228
rect 16836 27226 16892 27228
rect 16916 27226 16972 27228
rect 16996 27226 17052 27228
rect 16756 27174 16782 27226
rect 16782 27174 16812 27226
rect 16836 27174 16846 27226
rect 16846 27174 16892 27226
rect 16916 27174 16962 27226
rect 16962 27174 16972 27226
rect 16996 27174 17026 27226
rect 17026 27174 17052 27226
rect 16756 27172 16812 27174
rect 16836 27172 16892 27174
rect 16916 27172 16972 27174
rect 16996 27172 17052 27174
rect 19756 27226 19812 27228
rect 19836 27226 19892 27228
rect 19916 27226 19972 27228
rect 19996 27226 20052 27228
rect 19756 27174 19782 27226
rect 19782 27174 19812 27226
rect 19836 27174 19846 27226
rect 19846 27174 19892 27226
rect 19916 27174 19962 27226
rect 19962 27174 19972 27226
rect 19996 27174 20026 27226
rect 20026 27174 20052 27226
rect 19756 27172 19812 27174
rect 19836 27172 19892 27174
rect 19916 27172 19972 27174
rect 19996 27172 20052 27174
rect 3256 26682 3312 26684
rect 3336 26682 3392 26684
rect 3416 26682 3472 26684
rect 3496 26682 3552 26684
rect 3256 26630 3282 26682
rect 3282 26630 3312 26682
rect 3336 26630 3346 26682
rect 3346 26630 3392 26682
rect 3416 26630 3462 26682
rect 3462 26630 3472 26682
rect 3496 26630 3526 26682
rect 3526 26630 3552 26682
rect 3256 26628 3312 26630
rect 3336 26628 3392 26630
rect 3416 26628 3472 26630
rect 3496 26628 3552 26630
rect 6256 26682 6312 26684
rect 6336 26682 6392 26684
rect 6416 26682 6472 26684
rect 6496 26682 6552 26684
rect 6256 26630 6282 26682
rect 6282 26630 6312 26682
rect 6336 26630 6346 26682
rect 6346 26630 6392 26682
rect 6416 26630 6462 26682
rect 6462 26630 6472 26682
rect 6496 26630 6526 26682
rect 6526 26630 6552 26682
rect 6256 26628 6312 26630
rect 6336 26628 6392 26630
rect 6416 26628 6472 26630
rect 6496 26628 6552 26630
rect 9256 26682 9312 26684
rect 9336 26682 9392 26684
rect 9416 26682 9472 26684
rect 9496 26682 9552 26684
rect 9256 26630 9282 26682
rect 9282 26630 9312 26682
rect 9336 26630 9346 26682
rect 9346 26630 9392 26682
rect 9416 26630 9462 26682
rect 9462 26630 9472 26682
rect 9496 26630 9526 26682
rect 9526 26630 9552 26682
rect 9256 26628 9312 26630
rect 9336 26628 9392 26630
rect 9416 26628 9472 26630
rect 9496 26628 9552 26630
rect 12256 26682 12312 26684
rect 12336 26682 12392 26684
rect 12416 26682 12472 26684
rect 12496 26682 12552 26684
rect 12256 26630 12282 26682
rect 12282 26630 12312 26682
rect 12336 26630 12346 26682
rect 12346 26630 12392 26682
rect 12416 26630 12462 26682
rect 12462 26630 12472 26682
rect 12496 26630 12526 26682
rect 12526 26630 12552 26682
rect 12256 26628 12312 26630
rect 12336 26628 12392 26630
rect 12416 26628 12472 26630
rect 12496 26628 12552 26630
rect 15256 26682 15312 26684
rect 15336 26682 15392 26684
rect 15416 26682 15472 26684
rect 15496 26682 15552 26684
rect 15256 26630 15282 26682
rect 15282 26630 15312 26682
rect 15336 26630 15346 26682
rect 15346 26630 15392 26682
rect 15416 26630 15462 26682
rect 15462 26630 15472 26682
rect 15496 26630 15526 26682
rect 15526 26630 15552 26682
rect 15256 26628 15312 26630
rect 15336 26628 15392 26630
rect 15416 26628 15472 26630
rect 15496 26628 15552 26630
rect 18256 26682 18312 26684
rect 18336 26682 18392 26684
rect 18416 26682 18472 26684
rect 18496 26682 18552 26684
rect 18256 26630 18282 26682
rect 18282 26630 18312 26682
rect 18336 26630 18346 26682
rect 18346 26630 18392 26682
rect 18416 26630 18462 26682
rect 18462 26630 18472 26682
rect 18496 26630 18526 26682
rect 18526 26630 18552 26682
rect 18256 26628 18312 26630
rect 18336 26628 18392 26630
rect 18416 26628 18472 26630
rect 18496 26628 18552 26630
rect 21256 26682 21312 26684
rect 21336 26682 21392 26684
rect 21416 26682 21472 26684
rect 21496 26682 21552 26684
rect 21256 26630 21282 26682
rect 21282 26630 21312 26682
rect 21336 26630 21346 26682
rect 21346 26630 21392 26682
rect 21416 26630 21462 26682
rect 21462 26630 21472 26682
rect 21496 26630 21526 26682
rect 21526 26630 21552 26682
rect 21256 26628 21312 26630
rect 21336 26628 21392 26630
rect 21416 26628 21472 26630
rect 21496 26628 21552 26630
rect 1756 26138 1812 26140
rect 1836 26138 1892 26140
rect 1916 26138 1972 26140
rect 1996 26138 2052 26140
rect 1756 26086 1782 26138
rect 1782 26086 1812 26138
rect 1836 26086 1846 26138
rect 1846 26086 1892 26138
rect 1916 26086 1962 26138
rect 1962 26086 1972 26138
rect 1996 26086 2026 26138
rect 2026 26086 2052 26138
rect 1756 26084 1812 26086
rect 1836 26084 1892 26086
rect 1916 26084 1972 26086
rect 1996 26084 2052 26086
rect 4756 26138 4812 26140
rect 4836 26138 4892 26140
rect 4916 26138 4972 26140
rect 4996 26138 5052 26140
rect 4756 26086 4782 26138
rect 4782 26086 4812 26138
rect 4836 26086 4846 26138
rect 4846 26086 4892 26138
rect 4916 26086 4962 26138
rect 4962 26086 4972 26138
rect 4996 26086 5026 26138
rect 5026 26086 5052 26138
rect 4756 26084 4812 26086
rect 4836 26084 4892 26086
rect 4916 26084 4972 26086
rect 4996 26084 5052 26086
rect 7756 26138 7812 26140
rect 7836 26138 7892 26140
rect 7916 26138 7972 26140
rect 7996 26138 8052 26140
rect 7756 26086 7782 26138
rect 7782 26086 7812 26138
rect 7836 26086 7846 26138
rect 7846 26086 7892 26138
rect 7916 26086 7962 26138
rect 7962 26086 7972 26138
rect 7996 26086 8026 26138
rect 8026 26086 8052 26138
rect 7756 26084 7812 26086
rect 7836 26084 7892 26086
rect 7916 26084 7972 26086
rect 7996 26084 8052 26086
rect 10756 26138 10812 26140
rect 10836 26138 10892 26140
rect 10916 26138 10972 26140
rect 10996 26138 11052 26140
rect 10756 26086 10782 26138
rect 10782 26086 10812 26138
rect 10836 26086 10846 26138
rect 10846 26086 10892 26138
rect 10916 26086 10962 26138
rect 10962 26086 10972 26138
rect 10996 26086 11026 26138
rect 11026 26086 11052 26138
rect 10756 26084 10812 26086
rect 10836 26084 10892 26086
rect 10916 26084 10972 26086
rect 10996 26084 11052 26086
rect 13756 26138 13812 26140
rect 13836 26138 13892 26140
rect 13916 26138 13972 26140
rect 13996 26138 14052 26140
rect 13756 26086 13782 26138
rect 13782 26086 13812 26138
rect 13836 26086 13846 26138
rect 13846 26086 13892 26138
rect 13916 26086 13962 26138
rect 13962 26086 13972 26138
rect 13996 26086 14026 26138
rect 14026 26086 14052 26138
rect 13756 26084 13812 26086
rect 13836 26084 13892 26086
rect 13916 26084 13972 26086
rect 13996 26084 14052 26086
rect 16756 26138 16812 26140
rect 16836 26138 16892 26140
rect 16916 26138 16972 26140
rect 16996 26138 17052 26140
rect 16756 26086 16782 26138
rect 16782 26086 16812 26138
rect 16836 26086 16846 26138
rect 16846 26086 16892 26138
rect 16916 26086 16962 26138
rect 16962 26086 16972 26138
rect 16996 26086 17026 26138
rect 17026 26086 17052 26138
rect 16756 26084 16812 26086
rect 16836 26084 16892 26086
rect 16916 26084 16972 26086
rect 16996 26084 17052 26086
rect 19756 26138 19812 26140
rect 19836 26138 19892 26140
rect 19916 26138 19972 26140
rect 19996 26138 20052 26140
rect 19756 26086 19782 26138
rect 19782 26086 19812 26138
rect 19836 26086 19846 26138
rect 19846 26086 19892 26138
rect 19916 26086 19962 26138
rect 19962 26086 19972 26138
rect 19996 26086 20026 26138
rect 20026 26086 20052 26138
rect 19756 26084 19812 26086
rect 19836 26084 19892 26086
rect 19916 26084 19972 26086
rect 19996 26084 20052 26086
rect 3256 25594 3312 25596
rect 3336 25594 3392 25596
rect 3416 25594 3472 25596
rect 3496 25594 3552 25596
rect 3256 25542 3282 25594
rect 3282 25542 3312 25594
rect 3336 25542 3346 25594
rect 3346 25542 3392 25594
rect 3416 25542 3462 25594
rect 3462 25542 3472 25594
rect 3496 25542 3526 25594
rect 3526 25542 3552 25594
rect 3256 25540 3312 25542
rect 3336 25540 3392 25542
rect 3416 25540 3472 25542
rect 3496 25540 3552 25542
rect 6256 25594 6312 25596
rect 6336 25594 6392 25596
rect 6416 25594 6472 25596
rect 6496 25594 6552 25596
rect 6256 25542 6282 25594
rect 6282 25542 6312 25594
rect 6336 25542 6346 25594
rect 6346 25542 6392 25594
rect 6416 25542 6462 25594
rect 6462 25542 6472 25594
rect 6496 25542 6526 25594
rect 6526 25542 6552 25594
rect 6256 25540 6312 25542
rect 6336 25540 6392 25542
rect 6416 25540 6472 25542
rect 6496 25540 6552 25542
rect 9256 25594 9312 25596
rect 9336 25594 9392 25596
rect 9416 25594 9472 25596
rect 9496 25594 9552 25596
rect 9256 25542 9282 25594
rect 9282 25542 9312 25594
rect 9336 25542 9346 25594
rect 9346 25542 9392 25594
rect 9416 25542 9462 25594
rect 9462 25542 9472 25594
rect 9496 25542 9526 25594
rect 9526 25542 9552 25594
rect 9256 25540 9312 25542
rect 9336 25540 9392 25542
rect 9416 25540 9472 25542
rect 9496 25540 9552 25542
rect 12256 25594 12312 25596
rect 12336 25594 12392 25596
rect 12416 25594 12472 25596
rect 12496 25594 12552 25596
rect 12256 25542 12282 25594
rect 12282 25542 12312 25594
rect 12336 25542 12346 25594
rect 12346 25542 12392 25594
rect 12416 25542 12462 25594
rect 12462 25542 12472 25594
rect 12496 25542 12526 25594
rect 12526 25542 12552 25594
rect 12256 25540 12312 25542
rect 12336 25540 12392 25542
rect 12416 25540 12472 25542
rect 12496 25540 12552 25542
rect 15256 25594 15312 25596
rect 15336 25594 15392 25596
rect 15416 25594 15472 25596
rect 15496 25594 15552 25596
rect 15256 25542 15282 25594
rect 15282 25542 15312 25594
rect 15336 25542 15346 25594
rect 15346 25542 15392 25594
rect 15416 25542 15462 25594
rect 15462 25542 15472 25594
rect 15496 25542 15526 25594
rect 15526 25542 15552 25594
rect 15256 25540 15312 25542
rect 15336 25540 15392 25542
rect 15416 25540 15472 25542
rect 15496 25540 15552 25542
rect 18256 25594 18312 25596
rect 18336 25594 18392 25596
rect 18416 25594 18472 25596
rect 18496 25594 18552 25596
rect 18256 25542 18282 25594
rect 18282 25542 18312 25594
rect 18336 25542 18346 25594
rect 18346 25542 18392 25594
rect 18416 25542 18462 25594
rect 18462 25542 18472 25594
rect 18496 25542 18526 25594
rect 18526 25542 18552 25594
rect 18256 25540 18312 25542
rect 18336 25540 18392 25542
rect 18416 25540 18472 25542
rect 18496 25540 18552 25542
rect 21256 25594 21312 25596
rect 21336 25594 21392 25596
rect 21416 25594 21472 25596
rect 21496 25594 21552 25596
rect 21256 25542 21282 25594
rect 21282 25542 21312 25594
rect 21336 25542 21346 25594
rect 21346 25542 21392 25594
rect 21416 25542 21462 25594
rect 21462 25542 21472 25594
rect 21496 25542 21526 25594
rect 21526 25542 21552 25594
rect 21256 25540 21312 25542
rect 21336 25540 21392 25542
rect 21416 25540 21472 25542
rect 21496 25540 21552 25542
rect 1756 25050 1812 25052
rect 1836 25050 1892 25052
rect 1916 25050 1972 25052
rect 1996 25050 2052 25052
rect 1756 24998 1782 25050
rect 1782 24998 1812 25050
rect 1836 24998 1846 25050
rect 1846 24998 1892 25050
rect 1916 24998 1962 25050
rect 1962 24998 1972 25050
rect 1996 24998 2026 25050
rect 2026 24998 2052 25050
rect 1756 24996 1812 24998
rect 1836 24996 1892 24998
rect 1916 24996 1972 24998
rect 1996 24996 2052 24998
rect 4756 25050 4812 25052
rect 4836 25050 4892 25052
rect 4916 25050 4972 25052
rect 4996 25050 5052 25052
rect 4756 24998 4782 25050
rect 4782 24998 4812 25050
rect 4836 24998 4846 25050
rect 4846 24998 4892 25050
rect 4916 24998 4962 25050
rect 4962 24998 4972 25050
rect 4996 24998 5026 25050
rect 5026 24998 5052 25050
rect 4756 24996 4812 24998
rect 4836 24996 4892 24998
rect 4916 24996 4972 24998
rect 4996 24996 5052 24998
rect 7756 25050 7812 25052
rect 7836 25050 7892 25052
rect 7916 25050 7972 25052
rect 7996 25050 8052 25052
rect 7756 24998 7782 25050
rect 7782 24998 7812 25050
rect 7836 24998 7846 25050
rect 7846 24998 7892 25050
rect 7916 24998 7962 25050
rect 7962 24998 7972 25050
rect 7996 24998 8026 25050
rect 8026 24998 8052 25050
rect 7756 24996 7812 24998
rect 7836 24996 7892 24998
rect 7916 24996 7972 24998
rect 7996 24996 8052 24998
rect 10756 25050 10812 25052
rect 10836 25050 10892 25052
rect 10916 25050 10972 25052
rect 10996 25050 11052 25052
rect 10756 24998 10782 25050
rect 10782 24998 10812 25050
rect 10836 24998 10846 25050
rect 10846 24998 10892 25050
rect 10916 24998 10962 25050
rect 10962 24998 10972 25050
rect 10996 24998 11026 25050
rect 11026 24998 11052 25050
rect 10756 24996 10812 24998
rect 10836 24996 10892 24998
rect 10916 24996 10972 24998
rect 10996 24996 11052 24998
rect 13756 25050 13812 25052
rect 13836 25050 13892 25052
rect 13916 25050 13972 25052
rect 13996 25050 14052 25052
rect 13756 24998 13782 25050
rect 13782 24998 13812 25050
rect 13836 24998 13846 25050
rect 13846 24998 13892 25050
rect 13916 24998 13962 25050
rect 13962 24998 13972 25050
rect 13996 24998 14026 25050
rect 14026 24998 14052 25050
rect 13756 24996 13812 24998
rect 13836 24996 13892 24998
rect 13916 24996 13972 24998
rect 13996 24996 14052 24998
rect 16756 25050 16812 25052
rect 16836 25050 16892 25052
rect 16916 25050 16972 25052
rect 16996 25050 17052 25052
rect 16756 24998 16782 25050
rect 16782 24998 16812 25050
rect 16836 24998 16846 25050
rect 16846 24998 16892 25050
rect 16916 24998 16962 25050
rect 16962 24998 16972 25050
rect 16996 24998 17026 25050
rect 17026 24998 17052 25050
rect 16756 24996 16812 24998
rect 16836 24996 16892 24998
rect 16916 24996 16972 24998
rect 16996 24996 17052 24998
rect 19756 25050 19812 25052
rect 19836 25050 19892 25052
rect 19916 25050 19972 25052
rect 19996 25050 20052 25052
rect 19756 24998 19782 25050
rect 19782 24998 19812 25050
rect 19836 24998 19846 25050
rect 19846 24998 19892 25050
rect 19916 24998 19962 25050
rect 19962 24998 19972 25050
rect 19996 24998 20026 25050
rect 20026 24998 20052 25050
rect 19756 24996 19812 24998
rect 19836 24996 19892 24998
rect 19916 24996 19972 24998
rect 19996 24996 20052 24998
rect 3256 24506 3312 24508
rect 3336 24506 3392 24508
rect 3416 24506 3472 24508
rect 3496 24506 3552 24508
rect 3256 24454 3282 24506
rect 3282 24454 3312 24506
rect 3336 24454 3346 24506
rect 3346 24454 3392 24506
rect 3416 24454 3462 24506
rect 3462 24454 3472 24506
rect 3496 24454 3526 24506
rect 3526 24454 3552 24506
rect 3256 24452 3312 24454
rect 3336 24452 3392 24454
rect 3416 24452 3472 24454
rect 3496 24452 3552 24454
rect 6256 24506 6312 24508
rect 6336 24506 6392 24508
rect 6416 24506 6472 24508
rect 6496 24506 6552 24508
rect 6256 24454 6282 24506
rect 6282 24454 6312 24506
rect 6336 24454 6346 24506
rect 6346 24454 6392 24506
rect 6416 24454 6462 24506
rect 6462 24454 6472 24506
rect 6496 24454 6526 24506
rect 6526 24454 6552 24506
rect 6256 24452 6312 24454
rect 6336 24452 6392 24454
rect 6416 24452 6472 24454
rect 6496 24452 6552 24454
rect 9256 24506 9312 24508
rect 9336 24506 9392 24508
rect 9416 24506 9472 24508
rect 9496 24506 9552 24508
rect 9256 24454 9282 24506
rect 9282 24454 9312 24506
rect 9336 24454 9346 24506
rect 9346 24454 9392 24506
rect 9416 24454 9462 24506
rect 9462 24454 9472 24506
rect 9496 24454 9526 24506
rect 9526 24454 9552 24506
rect 9256 24452 9312 24454
rect 9336 24452 9392 24454
rect 9416 24452 9472 24454
rect 9496 24452 9552 24454
rect 12256 24506 12312 24508
rect 12336 24506 12392 24508
rect 12416 24506 12472 24508
rect 12496 24506 12552 24508
rect 12256 24454 12282 24506
rect 12282 24454 12312 24506
rect 12336 24454 12346 24506
rect 12346 24454 12392 24506
rect 12416 24454 12462 24506
rect 12462 24454 12472 24506
rect 12496 24454 12526 24506
rect 12526 24454 12552 24506
rect 12256 24452 12312 24454
rect 12336 24452 12392 24454
rect 12416 24452 12472 24454
rect 12496 24452 12552 24454
rect 15256 24506 15312 24508
rect 15336 24506 15392 24508
rect 15416 24506 15472 24508
rect 15496 24506 15552 24508
rect 15256 24454 15282 24506
rect 15282 24454 15312 24506
rect 15336 24454 15346 24506
rect 15346 24454 15392 24506
rect 15416 24454 15462 24506
rect 15462 24454 15472 24506
rect 15496 24454 15526 24506
rect 15526 24454 15552 24506
rect 15256 24452 15312 24454
rect 15336 24452 15392 24454
rect 15416 24452 15472 24454
rect 15496 24452 15552 24454
rect 18256 24506 18312 24508
rect 18336 24506 18392 24508
rect 18416 24506 18472 24508
rect 18496 24506 18552 24508
rect 18256 24454 18282 24506
rect 18282 24454 18312 24506
rect 18336 24454 18346 24506
rect 18346 24454 18392 24506
rect 18416 24454 18462 24506
rect 18462 24454 18472 24506
rect 18496 24454 18526 24506
rect 18526 24454 18552 24506
rect 18256 24452 18312 24454
rect 18336 24452 18392 24454
rect 18416 24452 18472 24454
rect 18496 24452 18552 24454
rect 21256 24506 21312 24508
rect 21336 24506 21392 24508
rect 21416 24506 21472 24508
rect 21496 24506 21552 24508
rect 21256 24454 21282 24506
rect 21282 24454 21312 24506
rect 21336 24454 21346 24506
rect 21346 24454 21392 24506
rect 21416 24454 21462 24506
rect 21462 24454 21472 24506
rect 21496 24454 21526 24506
rect 21526 24454 21552 24506
rect 21256 24452 21312 24454
rect 21336 24452 21392 24454
rect 21416 24452 21472 24454
rect 21496 24452 21552 24454
rect 1756 23962 1812 23964
rect 1836 23962 1892 23964
rect 1916 23962 1972 23964
rect 1996 23962 2052 23964
rect 1756 23910 1782 23962
rect 1782 23910 1812 23962
rect 1836 23910 1846 23962
rect 1846 23910 1892 23962
rect 1916 23910 1962 23962
rect 1962 23910 1972 23962
rect 1996 23910 2026 23962
rect 2026 23910 2052 23962
rect 1756 23908 1812 23910
rect 1836 23908 1892 23910
rect 1916 23908 1972 23910
rect 1996 23908 2052 23910
rect 4756 23962 4812 23964
rect 4836 23962 4892 23964
rect 4916 23962 4972 23964
rect 4996 23962 5052 23964
rect 4756 23910 4782 23962
rect 4782 23910 4812 23962
rect 4836 23910 4846 23962
rect 4846 23910 4892 23962
rect 4916 23910 4962 23962
rect 4962 23910 4972 23962
rect 4996 23910 5026 23962
rect 5026 23910 5052 23962
rect 4756 23908 4812 23910
rect 4836 23908 4892 23910
rect 4916 23908 4972 23910
rect 4996 23908 5052 23910
rect 7756 23962 7812 23964
rect 7836 23962 7892 23964
rect 7916 23962 7972 23964
rect 7996 23962 8052 23964
rect 7756 23910 7782 23962
rect 7782 23910 7812 23962
rect 7836 23910 7846 23962
rect 7846 23910 7892 23962
rect 7916 23910 7962 23962
rect 7962 23910 7972 23962
rect 7996 23910 8026 23962
rect 8026 23910 8052 23962
rect 7756 23908 7812 23910
rect 7836 23908 7892 23910
rect 7916 23908 7972 23910
rect 7996 23908 8052 23910
rect 10756 23962 10812 23964
rect 10836 23962 10892 23964
rect 10916 23962 10972 23964
rect 10996 23962 11052 23964
rect 10756 23910 10782 23962
rect 10782 23910 10812 23962
rect 10836 23910 10846 23962
rect 10846 23910 10892 23962
rect 10916 23910 10962 23962
rect 10962 23910 10972 23962
rect 10996 23910 11026 23962
rect 11026 23910 11052 23962
rect 10756 23908 10812 23910
rect 10836 23908 10892 23910
rect 10916 23908 10972 23910
rect 10996 23908 11052 23910
rect 13756 23962 13812 23964
rect 13836 23962 13892 23964
rect 13916 23962 13972 23964
rect 13996 23962 14052 23964
rect 13756 23910 13782 23962
rect 13782 23910 13812 23962
rect 13836 23910 13846 23962
rect 13846 23910 13892 23962
rect 13916 23910 13962 23962
rect 13962 23910 13972 23962
rect 13996 23910 14026 23962
rect 14026 23910 14052 23962
rect 13756 23908 13812 23910
rect 13836 23908 13892 23910
rect 13916 23908 13972 23910
rect 13996 23908 14052 23910
rect 16756 23962 16812 23964
rect 16836 23962 16892 23964
rect 16916 23962 16972 23964
rect 16996 23962 17052 23964
rect 16756 23910 16782 23962
rect 16782 23910 16812 23962
rect 16836 23910 16846 23962
rect 16846 23910 16892 23962
rect 16916 23910 16962 23962
rect 16962 23910 16972 23962
rect 16996 23910 17026 23962
rect 17026 23910 17052 23962
rect 16756 23908 16812 23910
rect 16836 23908 16892 23910
rect 16916 23908 16972 23910
rect 16996 23908 17052 23910
rect 19756 23962 19812 23964
rect 19836 23962 19892 23964
rect 19916 23962 19972 23964
rect 19996 23962 20052 23964
rect 19756 23910 19782 23962
rect 19782 23910 19812 23962
rect 19836 23910 19846 23962
rect 19846 23910 19892 23962
rect 19916 23910 19962 23962
rect 19962 23910 19972 23962
rect 19996 23910 20026 23962
rect 20026 23910 20052 23962
rect 19756 23908 19812 23910
rect 19836 23908 19892 23910
rect 19916 23908 19972 23910
rect 19996 23908 20052 23910
rect 3256 23418 3312 23420
rect 3336 23418 3392 23420
rect 3416 23418 3472 23420
rect 3496 23418 3552 23420
rect 3256 23366 3282 23418
rect 3282 23366 3312 23418
rect 3336 23366 3346 23418
rect 3346 23366 3392 23418
rect 3416 23366 3462 23418
rect 3462 23366 3472 23418
rect 3496 23366 3526 23418
rect 3526 23366 3552 23418
rect 3256 23364 3312 23366
rect 3336 23364 3392 23366
rect 3416 23364 3472 23366
rect 3496 23364 3552 23366
rect 6256 23418 6312 23420
rect 6336 23418 6392 23420
rect 6416 23418 6472 23420
rect 6496 23418 6552 23420
rect 6256 23366 6282 23418
rect 6282 23366 6312 23418
rect 6336 23366 6346 23418
rect 6346 23366 6392 23418
rect 6416 23366 6462 23418
rect 6462 23366 6472 23418
rect 6496 23366 6526 23418
rect 6526 23366 6552 23418
rect 6256 23364 6312 23366
rect 6336 23364 6392 23366
rect 6416 23364 6472 23366
rect 6496 23364 6552 23366
rect 9256 23418 9312 23420
rect 9336 23418 9392 23420
rect 9416 23418 9472 23420
rect 9496 23418 9552 23420
rect 9256 23366 9282 23418
rect 9282 23366 9312 23418
rect 9336 23366 9346 23418
rect 9346 23366 9392 23418
rect 9416 23366 9462 23418
rect 9462 23366 9472 23418
rect 9496 23366 9526 23418
rect 9526 23366 9552 23418
rect 9256 23364 9312 23366
rect 9336 23364 9392 23366
rect 9416 23364 9472 23366
rect 9496 23364 9552 23366
rect 12256 23418 12312 23420
rect 12336 23418 12392 23420
rect 12416 23418 12472 23420
rect 12496 23418 12552 23420
rect 12256 23366 12282 23418
rect 12282 23366 12312 23418
rect 12336 23366 12346 23418
rect 12346 23366 12392 23418
rect 12416 23366 12462 23418
rect 12462 23366 12472 23418
rect 12496 23366 12526 23418
rect 12526 23366 12552 23418
rect 12256 23364 12312 23366
rect 12336 23364 12392 23366
rect 12416 23364 12472 23366
rect 12496 23364 12552 23366
rect 15256 23418 15312 23420
rect 15336 23418 15392 23420
rect 15416 23418 15472 23420
rect 15496 23418 15552 23420
rect 15256 23366 15282 23418
rect 15282 23366 15312 23418
rect 15336 23366 15346 23418
rect 15346 23366 15392 23418
rect 15416 23366 15462 23418
rect 15462 23366 15472 23418
rect 15496 23366 15526 23418
rect 15526 23366 15552 23418
rect 15256 23364 15312 23366
rect 15336 23364 15392 23366
rect 15416 23364 15472 23366
rect 15496 23364 15552 23366
rect 18256 23418 18312 23420
rect 18336 23418 18392 23420
rect 18416 23418 18472 23420
rect 18496 23418 18552 23420
rect 18256 23366 18282 23418
rect 18282 23366 18312 23418
rect 18336 23366 18346 23418
rect 18346 23366 18392 23418
rect 18416 23366 18462 23418
rect 18462 23366 18472 23418
rect 18496 23366 18526 23418
rect 18526 23366 18552 23418
rect 18256 23364 18312 23366
rect 18336 23364 18392 23366
rect 18416 23364 18472 23366
rect 18496 23364 18552 23366
rect 21256 23418 21312 23420
rect 21336 23418 21392 23420
rect 21416 23418 21472 23420
rect 21496 23418 21552 23420
rect 21256 23366 21282 23418
rect 21282 23366 21312 23418
rect 21336 23366 21346 23418
rect 21346 23366 21392 23418
rect 21416 23366 21462 23418
rect 21462 23366 21472 23418
rect 21496 23366 21526 23418
rect 21526 23366 21552 23418
rect 21256 23364 21312 23366
rect 21336 23364 21392 23366
rect 21416 23364 21472 23366
rect 21496 23364 21552 23366
rect 1756 22874 1812 22876
rect 1836 22874 1892 22876
rect 1916 22874 1972 22876
rect 1996 22874 2052 22876
rect 1756 22822 1782 22874
rect 1782 22822 1812 22874
rect 1836 22822 1846 22874
rect 1846 22822 1892 22874
rect 1916 22822 1962 22874
rect 1962 22822 1972 22874
rect 1996 22822 2026 22874
rect 2026 22822 2052 22874
rect 1756 22820 1812 22822
rect 1836 22820 1892 22822
rect 1916 22820 1972 22822
rect 1996 22820 2052 22822
rect 4756 22874 4812 22876
rect 4836 22874 4892 22876
rect 4916 22874 4972 22876
rect 4996 22874 5052 22876
rect 4756 22822 4782 22874
rect 4782 22822 4812 22874
rect 4836 22822 4846 22874
rect 4846 22822 4892 22874
rect 4916 22822 4962 22874
rect 4962 22822 4972 22874
rect 4996 22822 5026 22874
rect 5026 22822 5052 22874
rect 4756 22820 4812 22822
rect 4836 22820 4892 22822
rect 4916 22820 4972 22822
rect 4996 22820 5052 22822
rect 7756 22874 7812 22876
rect 7836 22874 7892 22876
rect 7916 22874 7972 22876
rect 7996 22874 8052 22876
rect 7756 22822 7782 22874
rect 7782 22822 7812 22874
rect 7836 22822 7846 22874
rect 7846 22822 7892 22874
rect 7916 22822 7962 22874
rect 7962 22822 7972 22874
rect 7996 22822 8026 22874
rect 8026 22822 8052 22874
rect 7756 22820 7812 22822
rect 7836 22820 7892 22822
rect 7916 22820 7972 22822
rect 7996 22820 8052 22822
rect 10756 22874 10812 22876
rect 10836 22874 10892 22876
rect 10916 22874 10972 22876
rect 10996 22874 11052 22876
rect 10756 22822 10782 22874
rect 10782 22822 10812 22874
rect 10836 22822 10846 22874
rect 10846 22822 10892 22874
rect 10916 22822 10962 22874
rect 10962 22822 10972 22874
rect 10996 22822 11026 22874
rect 11026 22822 11052 22874
rect 10756 22820 10812 22822
rect 10836 22820 10892 22822
rect 10916 22820 10972 22822
rect 10996 22820 11052 22822
rect 13756 22874 13812 22876
rect 13836 22874 13892 22876
rect 13916 22874 13972 22876
rect 13996 22874 14052 22876
rect 13756 22822 13782 22874
rect 13782 22822 13812 22874
rect 13836 22822 13846 22874
rect 13846 22822 13892 22874
rect 13916 22822 13962 22874
rect 13962 22822 13972 22874
rect 13996 22822 14026 22874
rect 14026 22822 14052 22874
rect 13756 22820 13812 22822
rect 13836 22820 13892 22822
rect 13916 22820 13972 22822
rect 13996 22820 14052 22822
rect 16756 22874 16812 22876
rect 16836 22874 16892 22876
rect 16916 22874 16972 22876
rect 16996 22874 17052 22876
rect 16756 22822 16782 22874
rect 16782 22822 16812 22874
rect 16836 22822 16846 22874
rect 16846 22822 16892 22874
rect 16916 22822 16962 22874
rect 16962 22822 16972 22874
rect 16996 22822 17026 22874
rect 17026 22822 17052 22874
rect 16756 22820 16812 22822
rect 16836 22820 16892 22822
rect 16916 22820 16972 22822
rect 16996 22820 17052 22822
rect 19756 22874 19812 22876
rect 19836 22874 19892 22876
rect 19916 22874 19972 22876
rect 19996 22874 20052 22876
rect 19756 22822 19782 22874
rect 19782 22822 19812 22874
rect 19836 22822 19846 22874
rect 19846 22822 19892 22874
rect 19916 22822 19962 22874
rect 19962 22822 19972 22874
rect 19996 22822 20026 22874
rect 20026 22822 20052 22874
rect 19756 22820 19812 22822
rect 19836 22820 19892 22822
rect 19916 22820 19972 22822
rect 19996 22820 20052 22822
rect 3256 22330 3312 22332
rect 3336 22330 3392 22332
rect 3416 22330 3472 22332
rect 3496 22330 3552 22332
rect 3256 22278 3282 22330
rect 3282 22278 3312 22330
rect 3336 22278 3346 22330
rect 3346 22278 3392 22330
rect 3416 22278 3462 22330
rect 3462 22278 3472 22330
rect 3496 22278 3526 22330
rect 3526 22278 3552 22330
rect 3256 22276 3312 22278
rect 3336 22276 3392 22278
rect 3416 22276 3472 22278
rect 3496 22276 3552 22278
rect 6256 22330 6312 22332
rect 6336 22330 6392 22332
rect 6416 22330 6472 22332
rect 6496 22330 6552 22332
rect 6256 22278 6282 22330
rect 6282 22278 6312 22330
rect 6336 22278 6346 22330
rect 6346 22278 6392 22330
rect 6416 22278 6462 22330
rect 6462 22278 6472 22330
rect 6496 22278 6526 22330
rect 6526 22278 6552 22330
rect 6256 22276 6312 22278
rect 6336 22276 6392 22278
rect 6416 22276 6472 22278
rect 6496 22276 6552 22278
rect 9256 22330 9312 22332
rect 9336 22330 9392 22332
rect 9416 22330 9472 22332
rect 9496 22330 9552 22332
rect 9256 22278 9282 22330
rect 9282 22278 9312 22330
rect 9336 22278 9346 22330
rect 9346 22278 9392 22330
rect 9416 22278 9462 22330
rect 9462 22278 9472 22330
rect 9496 22278 9526 22330
rect 9526 22278 9552 22330
rect 9256 22276 9312 22278
rect 9336 22276 9392 22278
rect 9416 22276 9472 22278
rect 9496 22276 9552 22278
rect 12256 22330 12312 22332
rect 12336 22330 12392 22332
rect 12416 22330 12472 22332
rect 12496 22330 12552 22332
rect 12256 22278 12282 22330
rect 12282 22278 12312 22330
rect 12336 22278 12346 22330
rect 12346 22278 12392 22330
rect 12416 22278 12462 22330
rect 12462 22278 12472 22330
rect 12496 22278 12526 22330
rect 12526 22278 12552 22330
rect 12256 22276 12312 22278
rect 12336 22276 12392 22278
rect 12416 22276 12472 22278
rect 12496 22276 12552 22278
rect 15256 22330 15312 22332
rect 15336 22330 15392 22332
rect 15416 22330 15472 22332
rect 15496 22330 15552 22332
rect 15256 22278 15282 22330
rect 15282 22278 15312 22330
rect 15336 22278 15346 22330
rect 15346 22278 15392 22330
rect 15416 22278 15462 22330
rect 15462 22278 15472 22330
rect 15496 22278 15526 22330
rect 15526 22278 15552 22330
rect 15256 22276 15312 22278
rect 15336 22276 15392 22278
rect 15416 22276 15472 22278
rect 15496 22276 15552 22278
rect 18256 22330 18312 22332
rect 18336 22330 18392 22332
rect 18416 22330 18472 22332
rect 18496 22330 18552 22332
rect 18256 22278 18282 22330
rect 18282 22278 18312 22330
rect 18336 22278 18346 22330
rect 18346 22278 18392 22330
rect 18416 22278 18462 22330
rect 18462 22278 18472 22330
rect 18496 22278 18526 22330
rect 18526 22278 18552 22330
rect 18256 22276 18312 22278
rect 18336 22276 18392 22278
rect 18416 22276 18472 22278
rect 18496 22276 18552 22278
rect 21256 22330 21312 22332
rect 21336 22330 21392 22332
rect 21416 22330 21472 22332
rect 21496 22330 21552 22332
rect 21256 22278 21282 22330
rect 21282 22278 21312 22330
rect 21336 22278 21346 22330
rect 21346 22278 21392 22330
rect 21416 22278 21462 22330
rect 21462 22278 21472 22330
rect 21496 22278 21526 22330
rect 21526 22278 21552 22330
rect 21256 22276 21312 22278
rect 21336 22276 21392 22278
rect 21416 22276 21472 22278
rect 21496 22276 21552 22278
rect 1756 21786 1812 21788
rect 1836 21786 1892 21788
rect 1916 21786 1972 21788
rect 1996 21786 2052 21788
rect 1756 21734 1782 21786
rect 1782 21734 1812 21786
rect 1836 21734 1846 21786
rect 1846 21734 1892 21786
rect 1916 21734 1962 21786
rect 1962 21734 1972 21786
rect 1996 21734 2026 21786
rect 2026 21734 2052 21786
rect 1756 21732 1812 21734
rect 1836 21732 1892 21734
rect 1916 21732 1972 21734
rect 1996 21732 2052 21734
rect 4756 21786 4812 21788
rect 4836 21786 4892 21788
rect 4916 21786 4972 21788
rect 4996 21786 5052 21788
rect 4756 21734 4782 21786
rect 4782 21734 4812 21786
rect 4836 21734 4846 21786
rect 4846 21734 4892 21786
rect 4916 21734 4962 21786
rect 4962 21734 4972 21786
rect 4996 21734 5026 21786
rect 5026 21734 5052 21786
rect 4756 21732 4812 21734
rect 4836 21732 4892 21734
rect 4916 21732 4972 21734
rect 4996 21732 5052 21734
rect 7756 21786 7812 21788
rect 7836 21786 7892 21788
rect 7916 21786 7972 21788
rect 7996 21786 8052 21788
rect 7756 21734 7782 21786
rect 7782 21734 7812 21786
rect 7836 21734 7846 21786
rect 7846 21734 7892 21786
rect 7916 21734 7962 21786
rect 7962 21734 7972 21786
rect 7996 21734 8026 21786
rect 8026 21734 8052 21786
rect 7756 21732 7812 21734
rect 7836 21732 7892 21734
rect 7916 21732 7972 21734
rect 7996 21732 8052 21734
rect 10756 21786 10812 21788
rect 10836 21786 10892 21788
rect 10916 21786 10972 21788
rect 10996 21786 11052 21788
rect 10756 21734 10782 21786
rect 10782 21734 10812 21786
rect 10836 21734 10846 21786
rect 10846 21734 10892 21786
rect 10916 21734 10962 21786
rect 10962 21734 10972 21786
rect 10996 21734 11026 21786
rect 11026 21734 11052 21786
rect 10756 21732 10812 21734
rect 10836 21732 10892 21734
rect 10916 21732 10972 21734
rect 10996 21732 11052 21734
rect 13756 21786 13812 21788
rect 13836 21786 13892 21788
rect 13916 21786 13972 21788
rect 13996 21786 14052 21788
rect 13756 21734 13782 21786
rect 13782 21734 13812 21786
rect 13836 21734 13846 21786
rect 13846 21734 13892 21786
rect 13916 21734 13962 21786
rect 13962 21734 13972 21786
rect 13996 21734 14026 21786
rect 14026 21734 14052 21786
rect 13756 21732 13812 21734
rect 13836 21732 13892 21734
rect 13916 21732 13972 21734
rect 13996 21732 14052 21734
rect 16756 21786 16812 21788
rect 16836 21786 16892 21788
rect 16916 21786 16972 21788
rect 16996 21786 17052 21788
rect 16756 21734 16782 21786
rect 16782 21734 16812 21786
rect 16836 21734 16846 21786
rect 16846 21734 16892 21786
rect 16916 21734 16962 21786
rect 16962 21734 16972 21786
rect 16996 21734 17026 21786
rect 17026 21734 17052 21786
rect 16756 21732 16812 21734
rect 16836 21732 16892 21734
rect 16916 21732 16972 21734
rect 16996 21732 17052 21734
rect 19756 21786 19812 21788
rect 19836 21786 19892 21788
rect 19916 21786 19972 21788
rect 19996 21786 20052 21788
rect 19756 21734 19782 21786
rect 19782 21734 19812 21786
rect 19836 21734 19846 21786
rect 19846 21734 19892 21786
rect 19916 21734 19962 21786
rect 19962 21734 19972 21786
rect 19996 21734 20026 21786
rect 20026 21734 20052 21786
rect 19756 21732 19812 21734
rect 19836 21732 19892 21734
rect 19916 21732 19972 21734
rect 19996 21732 20052 21734
rect 3256 21242 3312 21244
rect 3336 21242 3392 21244
rect 3416 21242 3472 21244
rect 3496 21242 3552 21244
rect 3256 21190 3282 21242
rect 3282 21190 3312 21242
rect 3336 21190 3346 21242
rect 3346 21190 3392 21242
rect 3416 21190 3462 21242
rect 3462 21190 3472 21242
rect 3496 21190 3526 21242
rect 3526 21190 3552 21242
rect 3256 21188 3312 21190
rect 3336 21188 3392 21190
rect 3416 21188 3472 21190
rect 3496 21188 3552 21190
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6416 21242 6472 21244
rect 6496 21242 6552 21244
rect 6256 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6416 21190 6462 21242
rect 6462 21190 6472 21242
rect 6496 21190 6526 21242
rect 6526 21190 6552 21242
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 6416 21188 6472 21190
rect 6496 21188 6552 21190
rect 9256 21242 9312 21244
rect 9336 21242 9392 21244
rect 9416 21242 9472 21244
rect 9496 21242 9552 21244
rect 9256 21190 9282 21242
rect 9282 21190 9312 21242
rect 9336 21190 9346 21242
rect 9346 21190 9392 21242
rect 9416 21190 9462 21242
rect 9462 21190 9472 21242
rect 9496 21190 9526 21242
rect 9526 21190 9552 21242
rect 9256 21188 9312 21190
rect 9336 21188 9392 21190
rect 9416 21188 9472 21190
rect 9496 21188 9552 21190
rect 12256 21242 12312 21244
rect 12336 21242 12392 21244
rect 12416 21242 12472 21244
rect 12496 21242 12552 21244
rect 12256 21190 12282 21242
rect 12282 21190 12312 21242
rect 12336 21190 12346 21242
rect 12346 21190 12392 21242
rect 12416 21190 12462 21242
rect 12462 21190 12472 21242
rect 12496 21190 12526 21242
rect 12526 21190 12552 21242
rect 12256 21188 12312 21190
rect 12336 21188 12392 21190
rect 12416 21188 12472 21190
rect 12496 21188 12552 21190
rect 15256 21242 15312 21244
rect 15336 21242 15392 21244
rect 15416 21242 15472 21244
rect 15496 21242 15552 21244
rect 15256 21190 15282 21242
rect 15282 21190 15312 21242
rect 15336 21190 15346 21242
rect 15346 21190 15392 21242
rect 15416 21190 15462 21242
rect 15462 21190 15472 21242
rect 15496 21190 15526 21242
rect 15526 21190 15552 21242
rect 15256 21188 15312 21190
rect 15336 21188 15392 21190
rect 15416 21188 15472 21190
rect 15496 21188 15552 21190
rect 18256 21242 18312 21244
rect 18336 21242 18392 21244
rect 18416 21242 18472 21244
rect 18496 21242 18552 21244
rect 18256 21190 18282 21242
rect 18282 21190 18312 21242
rect 18336 21190 18346 21242
rect 18346 21190 18392 21242
rect 18416 21190 18462 21242
rect 18462 21190 18472 21242
rect 18496 21190 18526 21242
rect 18526 21190 18552 21242
rect 18256 21188 18312 21190
rect 18336 21188 18392 21190
rect 18416 21188 18472 21190
rect 18496 21188 18552 21190
rect 21256 21242 21312 21244
rect 21336 21242 21392 21244
rect 21416 21242 21472 21244
rect 21496 21242 21552 21244
rect 21256 21190 21282 21242
rect 21282 21190 21312 21242
rect 21336 21190 21346 21242
rect 21346 21190 21392 21242
rect 21416 21190 21462 21242
rect 21462 21190 21472 21242
rect 21496 21190 21526 21242
rect 21526 21190 21552 21242
rect 21256 21188 21312 21190
rect 21336 21188 21392 21190
rect 21416 21188 21472 21190
rect 21496 21188 21552 21190
rect 1756 20698 1812 20700
rect 1836 20698 1892 20700
rect 1916 20698 1972 20700
rect 1996 20698 2052 20700
rect 1756 20646 1782 20698
rect 1782 20646 1812 20698
rect 1836 20646 1846 20698
rect 1846 20646 1892 20698
rect 1916 20646 1962 20698
rect 1962 20646 1972 20698
rect 1996 20646 2026 20698
rect 2026 20646 2052 20698
rect 1756 20644 1812 20646
rect 1836 20644 1892 20646
rect 1916 20644 1972 20646
rect 1996 20644 2052 20646
rect 4756 20698 4812 20700
rect 4836 20698 4892 20700
rect 4916 20698 4972 20700
rect 4996 20698 5052 20700
rect 4756 20646 4782 20698
rect 4782 20646 4812 20698
rect 4836 20646 4846 20698
rect 4846 20646 4892 20698
rect 4916 20646 4962 20698
rect 4962 20646 4972 20698
rect 4996 20646 5026 20698
rect 5026 20646 5052 20698
rect 4756 20644 4812 20646
rect 4836 20644 4892 20646
rect 4916 20644 4972 20646
rect 4996 20644 5052 20646
rect 7756 20698 7812 20700
rect 7836 20698 7892 20700
rect 7916 20698 7972 20700
rect 7996 20698 8052 20700
rect 7756 20646 7782 20698
rect 7782 20646 7812 20698
rect 7836 20646 7846 20698
rect 7846 20646 7892 20698
rect 7916 20646 7962 20698
rect 7962 20646 7972 20698
rect 7996 20646 8026 20698
rect 8026 20646 8052 20698
rect 7756 20644 7812 20646
rect 7836 20644 7892 20646
rect 7916 20644 7972 20646
rect 7996 20644 8052 20646
rect 10756 20698 10812 20700
rect 10836 20698 10892 20700
rect 10916 20698 10972 20700
rect 10996 20698 11052 20700
rect 10756 20646 10782 20698
rect 10782 20646 10812 20698
rect 10836 20646 10846 20698
rect 10846 20646 10892 20698
rect 10916 20646 10962 20698
rect 10962 20646 10972 20698
rect 10996 20646 11026 20698
rect 11026 20646 11052 20698
rect 10756 20644 10812 20646
rect 10836 20644 10892 20646
rect 10916 20644 10972 20646
rect 10996 20644 11052 20646
rect 13756 20698 13812 20700
rect 13836 20698 13892 20700
rect 13916 20698 13972 20700
rect 13996 20698 14052 20700
rect 13756 20646 13782 20698
rect 13782 20646 13812 20698
rect 13836 20646 13846 20698
rect 13846 20646 13892 20698
rect 13916 20646 13962 20698
rect 13962 20646 13972 20698
rect 13996 20646 14026 20698
rect 14026 20646 14052 20698
rect 13756 20644 13812 20646
rect 13836 20644 13892 20646
rect 13916 20644 13972 20646
rect 13996 20644 14052 20646
rect 16756 20698 16812 20700
rect 16836 20698 16892 20700
rect 16916 20698 16972 20700
rect 16996 20698 17052 20700
rect 16756 20646 16782 20698
rect 16782 20646 16812 20698
rect 16836 20646 16846 20698
rect 16846 20646 16892 20698
rect 16916 20646 16962 20698
rect 16962 20646 16972 20698
rect 16996 20646 17026 20698
rect 17026 20646 17052 20698
rect 16756 20644 16812 20646
rect 16836 20644 16892 20646
rect 16916 20644 16972 20646
rect 16996 20644 17052 20646
rect 19756 20698 19812 20700
rect 19836 20698 19892 20700
rect 19916 20698 19972 20700
rect 19996 20698 20052 20700
rect 19756 20646 19782 20698
rect 19782 20646 19812 20698
rect 19836 20646 19846 20698
rect 19846 20646 19892 20698
rect 19916 20646 19962 20698
rect 19962 20646 19972 20698
rect 19996 20646 20026 20698
rect 20026 20646 20052 20698
rect 19756 20644 19812 20646
rect 19836 20644 19892 20646
rect 19916 20644 19972 20646
rect 19996 20644 20052 20646
rect 3256 20154 3312 20156
rect 3336 20154 3392 20156
rect 3416 20154 3472 20156
rect 3496 20154 3552 20156
rect 3256 20102 3282 20154
rect 3282 20102 3312 20154
rect 3336 20102 3346 20154
rect 3346 20102 3392 20154
rect 3416 20102 3462 20154
rect 3462 20102 3472 20154
rect 3496 20102 3526 20154
rect 3526 20102 3552 20154
rect 3256 20100 3312 20102
rect 3336 20100 3392 20102
rect 3416 20100 3472 20102
rect 3496 20100 3552 20102
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6416 20154 6472 20156
rect 6496 20154 6552 20156
rect 6256 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6416 20102 6462 20154
rect 6462 20102 6472 20154
rect 6496 20102 6526 20154
rect 6526 20102 6552 20154
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 6416 20100 6472 20102
rect 6496 20100 6552 20102
rect 9256 20154 9312 20156
rect 9336 20154 9392 20156
rect 9416 20154 9472 20156
rect 9496 20154 9552 20156
rect 9256 20102 9282 20154
rect 9282 20102 9312 20154
rect 9336 20102 9346 20154
rect 9346 20102 9392 20154
rect 9416 20102 9462 20154
rect 9462 20102 9472 20154
rect 9496 20102 9526 20154
rect 9526 20102 9552 20154
rect 9256 20100 9312 20102
rect 9336 20100 9392 20102
rect 9416 20100 9472 20102
rect 9496 20100 9552 20102
rect 12256 20154 12312 20156
rect 12336 20154 12392 20156
rect 12416 20154 12472 20156
rect 12496 20154 12552 20156
rect 12256 20102 12282 20154
rect 12282 20102 12312 20154
rect 12336 20102 12346 20154
rect 12346 20102 12392 20154
rect 12416 20102 12462 20154
rect 12462 20102 12472 20154
rect 12496 20102 12526 20154
rect 12526 20102 12552 20154
rect 12256 20100 12312 20102
rect 12336 20100 12392 20102
rect 12416 20100 12472 20102
rect 12496 20100 12552 20102
rect 15256 20154 15312 20156
rect 15336 20154 15392 20156
rect 15416 20154 15472 20156
rect 15496 20154 15552 20156
rect 15256 20102 15282 20154
rect 15282 20102 15312 20154
rect 15336 20102 15346 20154
rect 15346 20102 15392 20154
rect 15416 20102 15462 20154
rect 15462 20102 15472 20154
rect 15496 20102 15526 20154
rect 15526 20102 15552 20154
rect 15256 20100 15312 20102
rect 15336 20100 15392 20102
rect 15416 20100 15472 20102
rect 15496 20100 15552 20102
rect 18256 20154 18312 20156
rect 18336 20154 18392 20156
rect 18416 20154 18472 20156
rect 18496 20154 18552 20156
rect 18256 20102 18282 20154
rect 18282 20102 18312 20154
rect 18336 20102 18346 20154
rect 18346 20102 18392 20154
rect 18416 20102 18462 20154
rect 18462 20102 18472 20154
rect 18496 20102 18526 20154
rect 18526 20102 18552 20154
rect 18256 20100 18312 20102
rect 18336 20100 18392 20102
rect 18416 20100 18472 20102
rect 18496 20100 18552 20102
rect 21256 20154 21312 20156
rect 21336 20154 21392 20156
rect 21416 20154 21472 20156
rect 21496 20154 21552 20156
rect 21256 20102 21282 20154
rect 21282 20102 21312 20154
rect 21336 20102 21346 20154
rect 21346 20102 21392 20154
rect 21416 20102 21462 20154
rect 21462 20102 21472 20154
rect 21496 20102 21526 20154
rect 21526 20102 21552 20154
rect 21256 20100 21312 20102
rect 21336 20100 21392 20102
rect 21416 20100 21472 20102
rect 21496 20100 21552 20102
rect 1756 19610 1812 19612
rect 1836 19610 1892 19612
rect 1916 19610 1972 19612
rect 1996 19610 2052 19612
rect 1756 19558 1782 19610
rect 1782 19558 1812 19610
rect 1836 19558 1846 19610
rect 1846 19558 1892 19610
rect 1916 19558 1962 19610
rect 1962 19558 1972 19610
rect 1996 19558 2026 19610
rect 2026 19558 2052 19610
rect 1756 19556 1812 19558
rect 1836 19556 1892 19558
rect 1916 19556 1972 19558
rect 1996 19556 2052 19558
rect 4756 19610 4812 19612
rect 4836 19610 4892 19612
rect 4916 19610 4972 19612
rect 4996 19610 5052 19612
rect 4756 19558 4782 19610
rect 4782 19558 4812 19610
rect 4836 19558 4846 19610
rect 4846 19558 4892 19610
rect 4916 19558 4962 19610
rect 4962 19558 4972 19610
rect 4996 19558 5026 19610
rect 5026 19558 5052 19610
rect 4756 19556 4812 19558
rect 4836 19556 4892 19558
rect 4916 19556 4972 19558
rect 4996 19556 5052 19558
rect 7756 19610 7812 19612
rect 7836 19610 7892 19612
rect 7916 19610 7972 19612
rect 7996 19610 8052 19612
rect 7756 19558 7782 19610
rect 7782 19558 7812 19610
rect 7836 19558 7846 19610
rect 7846 19558 7892 19610
rect 7916 19558 7962 19610
rect 7962 19558 7972 19610
rect 7996 19558 8026 19610
rect 8026 19558 8052 19610
rect 7756 19556 7812 19558
rect 7836 19556 7892 19558
rect 7916 19556 7972 19558
rect 7996 19556 8052 19558
rect 10756 19610 10812 19612
rect 10836 19610 10892 19612
rect 10916 19610 10972 19612
rect 10996 19610 11052 19612
rect 10756 19558 10782 19610
rect 10782 19558 10812 19610
rect 10836 19558 10846 19610
rect 10846 19558 10892 19610
rect 10916 19558 10962 19610
rect 10962 19558 10972 19610
rect 10996 19558 11026 19610
rect 11026 19558 11052 19610
rect 10756 19556 10812 19558
rect 10836 19556 10892 19558
rect 10916 19556 10972 19558
rect 10996 19556 11052 19558
rect 13756 19610 13812 19612
rect 13836 19610 13892 19612
rect 13916 19610 13972 19612
rect 13996 19610 14052 19612
rect 13756 19558 13782 19610
rect 13782 19558 13812 19610
rect 13836 19558 13846 19610
rect 13846 19558 13892 19610
rect 13916 19558 13962 19610
rect 13962 19558 13972 19610
rect 13996 19558 14026 19610
rect 14026 19558 14052 19610
rect 13756 19556 13812 19558
rect 13836 19556 13892 19558
rect 13916 19556 13972 19558
rect 13996 19556 14052 19558
rect 16756 19610 16812 19612
rect 16836 19610 16892 19612
rect 16916 19610 16972 19612
rect 16996 19610 17052 19612
rect 16756 19558 16782 19610
rect 16782 19558 16812 19610
rect 16836 19558 16846 19610
rect 16846 19558 16892 19610
rect 16916 19558 16962 19610
rect 16962 19558 16972 19610
rect 16996 19558 17026 19610
rect 17026 19558 17052 19610
rect 16756 19556 16812 19558
rect 16836 19556 16892 19558
rect 16916 19556 16972 19558
rect 16996 19556 17052 19558
rect 19756 19610 19812 19612
rect 19836 19610 19892 19612
rect 19916 19610 19972 19612
rect 19996 19610 20052 19612
rect 19756 19558 19782 19610
rect 19782 19558 19812 19610
rect 19836 19558 19846 19610
rect 19846 19558 19892 19610
rect 19916 19558 19962 19610
rect 19962 19558 19972 19610
rect 19996 19558 20026 19610
rect 20026 19558 20052 19610
rect 19756 19556 19812 19558
rect 19836 19556 19892 19558
rect 19916 19556 19972 19558
rect 19996 19556 20052 19558
rect 3256 19066 3312 19068
rect 3336 19066 3392 19068
rect 3416 19066 3472 19068
rect 3496 19066 3552 19068
rect 3256 19014 3282 19066
rect 3282 19014 3312 19066
rect 3336 19014 3346 19066
rect 3346 19014 3392 19066
rect 3416 19014 3462 19066
rect 3462 19014 3472 19066
rect 3496 19014 3526 19066
rect 3526 19014 3552 19066
rect 3256 19012 3312 19014
rect 3336 19012 3392 19014
rect 3416 19012 3472 19014
rect 3496 19012 3552 19014
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6416 19066 6472 19068
rect 6496 19066 6552 19068
rect 6256 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6416 19014 6462 19066
rect 6462 19014 6472 19066
rect 6496 19014 6526 19066
rect 6526 19014 6552 19066
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 6416 19012 6472 19014
rect 6496 19012 6552 19014
rect 9256 19066 9312 19068
rect 9336 19066 9392 19068
rect 9416 19066 9472 19068
rect 9496 19066 9552 19068
rect 9256 19014 9282 19066
rect 9282 19014 9312 19066
rect 9336 19014 9346 19066
rect 9346 19014 9392 19066
rect 9416 19014 9462 19066
rect 9462 19014 9472 19066
rect 9496 19014 9526 19066
rect 9526 19014 9552 19066
rect 9256 19012 9312 19014
rect 9336 19012 9392 19014
rect 9416 19012 9472 19014
rect 9496 19012 9552 19014
rect 12256 19066 12312 19068
rect 12336 19066 12392 19068
rect 12416 19066 12472 19068
rect 12496 19066 12552 19068
rect 12256 19014 12282 19066
rect 12282 19014 12312 19066
rect 12336 19014 12346 19066
rect 12346 19014 12392 19066
rect 12416 19014 12462 19066
rect 12462 19014 12472 19066
rect 12496 19014 12526 19066
rect 12526 19014 12552 19066
rect 12256 19012 12312 19014
rect 12336 19012 12392 19014
rect 12416 19012 12472 19014
rect 12496 19012 12552 19014
rect 15256 19066 15312 19068
rect 15336 19066 15392 19068
rect 15416 19066 15472 19068
rect 15496 19066 15552 19068
rect 15256 19014 15282 19066
rect 15282 19014 15312 19066
rect 15336 19014 15346 19066
rect 15346 19014 15392 19066
rect 15416 19014 15462 19066
rect 15462 19014 15472 19066
rect 15496 19014 15526 19066
rect 15526 19014 15552 19066
rect 15256 19012 15312 19014
rect 15336 19012 15392 19014
rect 15416 19012 15472 19014
rect 15496 19012 15552 19014
rect 18256 19066 18312 19068
rect 18336 19066 18392 19068
rect 18416 19066 18472 19068
rect 18496 19066 18552 19068
rect 18256 19014 18282 19066
rect 18282 19014 18312 19066
rect 18336 19014 18346 19066
rect 18346 19014 18392 19066
rect 18416 19014 18462 19066
rect 18462 19014 18472 19066
rect 18496 19014 18526 19066
rect 18526 19014 18552 19066
rect 18256 19012 18312 19014
rect 18336 19012 18392 19014
rect 18416 19012 18472 19014
rect 18496 19012 18552 19014
rect 21256 19066 21312 19068
rect 21336 19066 21392 19068
rect 21416 19066 21472 19068
rect 21496 19066 21552 19068
rect 21256 19014 21282 19066
rect 21282 19014 21312 19066
rect 21336 19014 21346 19066
rect 21346 19014 21392 19066
rect 21416 19014 21462 19066
rect 21462 19014 21472 19066
rect 21496 19014 21526 19066
rect 21526 19014 21552 19066
rect 21256 19012 21312 19014
rect 21336 19012 21392 19014
rect 21416 19012 21472 19014
rect 21496 19012 21552 19014
rect 1756 18522 1812 18524
rect 1836 18522 1892 18524
rect 1916 18522 1972 18524
rect 1996 18522 2052 18524
rect 1756 18470 1782 18522
rect 1782 18470 1812 18522
rect 1836 18470 1846 18522
rect 1846 18470 1892 18522
rect 1916 18470 1962 18522
rect 1962 18470 1972 18522
rect 1996 18470 2026 18522
rect 2026 18470 2052 18522
rect 1756 18468 1812 18470
rect 1836 18468 1892 18470
rect 1916 18468 1972 18470
rect 1996 18468 2052 18470
rect 4756 18522 4812 18524
rect 4836 18522 4892 18524
rect 4916 18522 4972 18524
rect 4996 18522 5052 18524
rect 4756 18470 4782 18522
rect 4782 18470 4812 18522
rect 4836 18470 4846 18522
rect 4846 18470 4892 18522
rect 4916 18470 4962 18522
rect 4962 18470 4972 18522
rect 4996 18470 5026 18522
rect 5026 18470 5052 18522
rect 4756 18468 4812 18470
rect 4836 18468 4892 18470
rect 4916 18468 4972 18470
rect 4996 18468 5052 18470
rect 7756 18522 7812 18524
rect 7836 18522 7892 18524
rect 7916 18522 7972 18524
rect 7996 18522 8052 18524
rect 7756 18470 7782 18522
rect 7782 18470 7812 18522
rect 7836 18470 7846 18522
rect 7846 18470 7892 18522
rect 7916 18470 7962 18522
rect 7962 18470 7972 18522
rect 7996 18470 8026 18522
rect 8026 18470 8052 18522
rect 7756 18468 7812 18470
rect 7836 18468 7892 18470
rect 7916 18468 7972 18470
rect 7996 18468 8052 18470
rect 10756 18522 10812 18524
rect 10836 18522 10892 18524
rect 10916 18522 10972 18524
rect 10996 18522 11052 18524
rect 10756 18470 10782 18522
rect 10782 18470 10812 18522
rect 10836 18470 10846 18522
rect 10846 18470 10892 18522
rect 10916 18470 10962 18522
rect 10962 18470 10972 18522
rect 10996 18470 11026 18522
rect 11026 18470 11052 18522
rect 10756 18468 10812 18470
rect 10836 18468 10892 18470
rect 10916 18468 10972 18470
rect 10996 18468 11052 18470
rect 13756 18522 13812 18524
rect 13836 18522 13892 18524
rect 13916 18522 13972 18524
rect 13996 18522 14052 18524
rect 13756 18470 13782 18522
rect 13782 18470 13812 18522
rect 13836 18470 13846 18522
rect 13846 18470 13892 18522
rect 13916 18470 13962 18522
rect 13962 18470 13972 18522
rect 13996 18470 14026 18522
rect 14026 18470 14052 18522
rect 13756 18468 13812 18470
rect 13836 18468 13892 18470
rect 13916 18468 13972 18470
rect 13996 18468 14052 18470
rect 16756 18522 16812 18524
rect 16836 18522 16892 18524
rect 16916 18522 16972 18524
rect 16996 18522 17052 18524
rect 16756 18470 16782 18522
rect 16782 18470 16812 18522
rect 16836 18470 16846 18522
rect 16846 18470 16892 18522
rect 16916 18470 16962 18522
rect 16962 18470 16972 18522
rect 16996 18470 17026 18522
rect 17026 18470 17052 18522
rect 16756 18468 16812 18470
rect 16836 18468 16892 18470
rect 16916 18468 16972 18470
rect 16996 18468 17052 18470
rect 19756 18522 19812 18524
rect 19836 18522 19892 18524
rect 19916 18522 19972 18524
rect 19996 18522 20052 18524
rect 19756 18470 19782 18522
rect 19782 18470 19812 18522
rect 19836 18470 19846 18522
rect 19846 18470 19892 18522
rect 19916 18470 19962 18522
rect 19962 18470 19972 18522
rect 19996 18470 20026 18522
rect 20026 18470 20052 18522
rect 19756 18468 19812 18470
rect 19836 18468 19892 18470
rect 19916 18468 19972 18470
rect 19996 18468 20052 18470
rect 3256 17978 3312 17980
rect 3336 17978 3392 17980
rect 3416 17978 3472 17980
rect 3496 17978 3552 17980
rect 3256 17926 3282 17978
rect 3282 17926 3312 17978
rect 3336 17926 3346 17978
rect 3346 17926 3392 17978
rect 3416 17926 3462 17978
rect 3462 17926 3472 17978
rect 3496 17926 3526 17978
rect 3526 17926 3552 17978
rect 3256 17924 3312 17926
rect 3336 17924 3392 17926
rect 3416 17924 3472 17926
rect 3496 17924 3552 17926
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6416 17978 6472 17980
rect 6496 17978 6552 17980
rect 6256 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6416 17926 6462 17978
rect 6462 17926 6472 17978
rect 6496 17926 6526 17978
rect 6526 17926 6552 17978
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 6416 17924 6472 17926
rect 6496 17924 6552 17926
rect 9256 17978 9312 17980
rect 9336 17978 9392 17980
rect 9416 17978 9472 17980
rect 9496 17978 9552 17980
rect 9256 17926 9282 17978
rect 9282 17926 9312 17978
rect 9336 17926 9346 17978
rect 9346 17926 9392 17978
rect 9416 17926 9462 17978
rect 9462 17926 9472 17978
rect 9496 17926 9526 17978
rect 9526 17926 9552 17978
rect 9256 17924 9312 17926
rect 9336 17924 9392 17926
rect 9416 17924 9472 17926
rect 9496 17924 9552 17926
rect 12256 17978 12312 17980
rect 12336 17978 12392 17980
rect 12416 17978 12472 17980
rect 12496 17978 12552 17980
rect 12256 17926 12282 17978
rect 12282 17926 12312 17978
rect 12336 17926 12346 17978
rect 12346 17926 12392 17978
rect 12416 17926 12462 17978
rect 12462 17926 12472 17978
rect 12496 17926 12526 17978
rect 12526 17926 12552 17978
rect 12256 17924 12312 17926
rect 12336 17924 12392 17926
rect 12416 17924 12472 17926
rect 12496 17924 12552 17926
rect 15256 17978 15312 17980
rect 15336 17978 15392 17980
rect 15416 17978 15472 17980
rect 15496 17978 15552 17980
rect 15256 17926 15282 17978
rect 15282 17926 15312 17978
rect 15336 17926 15346 17978
rect 15346 17926 15392 17978
rect 15416 17926 15462 17978
rect 15462 17926 15472 17978
rect 15496 17926 15526 17978
rect 15526 17926 15552 17978
rect 15256 17924 15312 17926
rect 15336 17924 15392 17926
rect 15416 17924 15472 17926
rect 15496 17924 15552 17926
rect 18256 17978 18312 17980
rect 18336 17978 18392 17980
rect 18416 17978 18472 17980
rect 18496 17978 18552 17980
rect 18256 17926 18282 17978
rect 18282 17926 18312 17978
rect 18336 17926 18346 17978
rect 18346 17926 18392 17978
rect 18416 17926 18462 17978
rect 18462 17926 18472 17978
rect 18496 17926 18526 17978
rect 18526 17926 18552 17978
rect 18256 17924 18312 17926
rect 18336 17924 18392 17926
rect 18416 17924 18472 17926
rect 18496 17924 18552 17926
rect 21256 17978 21312 17980
rect 21336 17978 21392 17980
rect 21416 17978 21472 17980
rect 21496 17978 21552 17980
rect 21256 17926 21282 17978
rect 21282 17926 21312 17978
rect 21336 17926 21346 17978
rect 21346 17926 21392 17978
rect 21416 17926 21462 17978
rect 21462 17926 21472 17978
rect 21496 17926 21526 17978
rect 21526 17926 21552 17978
rect 21256 17924 21312 17926
rect 21336 17924 21392 17926
rect 21416 17924 21472 17926
rect 21496 17924 21552 17926
rect 1756 17434 1812 17436
rect 1836 17434 1892 17436
rect 1916 17434 1972 17436
rect 1996 17434 2052 17436
rect 1756 17382 1782 17434
rect 1782 17382 1812 17434
rect 1836 17382 1846 17434
rect 1846 17382 1892 17434
rect 1916 17382 1962 17434
rect 1962 17382 1972 17434
rect 1996 17382 2026 17434
rect 2026 17382 2052 17434
rect 1756 17380 1812 17382
rect 1836 17380 1892 17382
rect 1916 17380 1972 17382
rect 1996 17380 2052 17382
rect 4756 17434 4812 17436
rect 4836 17434 4892 17436
rect 4916 17434 4972 17436
rect 4996 17434 5052 17436
rect 4756 17382 4782 17434
rect 4782 17382 4812 17434
rect 4836 17382 4846 17434
rect 4846 17382 4892 17434
rect 4916 17382 4962 17434
rect 4962 17382 4972 17434
rect 4996 17382 5026 17434
rect 5026 17382 5052 17434
rect 4756 17380 4812 17382
rect 4836 17380 4892 17382
rect 4916 17380 4972 17382
rect 4996 17380 5052 17382
rect 7756 17434 7812 17436
rect 7836 17434 7892 17436
rect 7916 17434 7972 17436
rect 7996 17434 8052 17436
rect 7756 17382 7782 17434
rect 7782 17382 7812 17434
rect 7836 17382 7846 17434
rect 7846 17382 7892 17434
rect 7916 17382 7962 17434
rect 7962 17382 7972 17434
rect 7996 17382 8026 17434
rect 8026 17382 8052 17434
rect 7756 17380 7812 17382
rect 7836 17380 7892 17382
rect 7916 17380 7972 17382
rect 7996 17380 8052 17382
rect 10756 17434 10812 17436
rect 10836 17434 10892 17436
rect 10916 17434 10972 17436
rect 10996 17434 11052 17436
rect 10756 17382 10782 17434
rect 10782 17382 10812 17434
rect 10836 17382 10846 17434
rect 10846 17382 10892 17434
rect 10916 17382 10962 17434
rect 10962 17382 10972 17434
rect 10996 17382 11026 17434
rect 11026 17382 11052 17434
rect 10756 17380 10812 17382
rect 10836 17380 10892 17382
rect 10916 17380 10972 17382
rect 10996 17380 11052 17382
rect 13756 17434 13812 17436
rect 13836 17434 13892 17436
rect 13916 17434 13972 17436
rect 13996 17434 14052 17436
rect 13756 17382 13782 17434
rect 13782 17382 13812 17434
rect 13836 17382 13846 17434
rect 13846 17382 13892 17434
rect 13916 17382 13962 17434
rect 13962 17382 13972 17434
rect 13996 17382 14026 17434
rect 14026 17382 14052 17434
rect 13756 17380 13812 17382
rect 13836 17380 13892 17382
rect 13916 17380 13972 17382
rect 13996 17380 14052 17382
rect 16756 17434 16812 17436
rect 16836 17434 16892 17436
rect 16916 17434 16972 17436
rect 16996 17434 17052 17436
rect 16756 17382 16782 17434
rect 16782 17382 16812 17434
rect 16836 17382 16846 17434
rect 16846 17382 16892 17434
rect 16916 17382 16962 17434
rect 16962 17382 16972 17434
rect 16996 17382 17026 17434
rect 17026 17382 17052 17434
rect 16756 17380 16812 17382
rect 16836 17380 16892 17382
rect 16916 17380 16972 17382
rect 16996 17380 17052 17382
rect 19756 17434 19812 17436
rect 19836 17434 19892 17436
rect 19916 17434 19972 17436
rect 19996 17434 20052 17436
rect 19756 17382 19782 17434
rect 19782 17382 19812 17434
rect 19836 17382 19846 17434
rect 19846 17382 19892 17434
rect 19916 17382 19962 17434
rect 19962 17382 19972 17434
rect 19996 17382 20026 17434
rect 20026 17382 20052 17434
rect 19756 17380 19812 17382
rect 19836 17380 19892 17382
rect 19916 17380 19972 17382
rect 19996 17380 20052 17382
rect 3256 16890 3312 16892
rect 3336 16890 3392 16892
rect 3416 16890 3472 16892
rect 3496 16890 3552 16892
rect 3256 16838 3282 16890
rect 3282 16838 3312 16890
rect 3336 16838 3346 16890
rect 3346 16838 3392 16890
rect 3416 16838 3462 16890
rect 3462 16838 3472 16890
rect 3496 16838 3526 16890
rect 3526 16838 3552 16890
rect 3256 16836 3312 16838
rect 3336 16836 3392 16838
rect 3416 16836 3472 16838
rect 3496 16836 3552 16838
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6416 16890 6472 16892
rect 6496 16890 6552 16892
rect 6256 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6416 16838 6462 16890
rect 6462 16838 6472 16890
rect 6496 16838 6526 16890
rect 6526 16838 6552 16890
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6416 16836 6472 16838
rect 6496 16836 6552 16838
rect 9256 16890 9312 16892
rect 9336 16890 9392 16892
rect 9416 16890 9472 16892
rect 9496 16890 9552 16892
rect 9256 16838 9282 16890
rect 9282 16838 9312 16890
rect 9336 16838 9346 16890
rect 9346 16838 9392 16890
rect 9416 16838 9462 16890
rect 9462 16838 9472 16890
rect 9496 16838 9526 16890
rect 9526 16838 9552 16890
rect 9256 16836 9312 16838
rect 9336 16836 9392 16838
rect 9416 16836 9472 16838
rect 9496 16836 9552 16838
rect 12256 16890 12312 16892
rect 12336 16890 12392 16892
rect 12416 16890 12472 16892
rect 12496 16890 12552 16892
rect 12256 16838 12282 16890
rect 12282 16838 12312 16890
rect 12336 16838 12346 16890
rect 12346 16838 12392 16890
rect 12416 16838 12462 16890
rect 12462 16838 12472 16890
rect 12496 16838 12526 16890
rect 12526 16838 12552 16890
rect 12256 16836 12312 16838
rect 12336 16836 12392 16838
rect 12416 16836 12472 16838
rect 12496 16836 12552 16838
rect 15256 16890 15312 16892
rect 15336 16890 15392 16892
rect 15416 16890 15472 16892
rect 15496 16890 15552 16892
rect 15256 16838 15282 16890
rect 15282 16838 15312 16890
rect 15336 16838 15346 16890
rect 15346 16838 15392 16890
rect 15416 16838 15462 16890
rect 15462 16838 15472 16890
rect 15496 16838 15526 16890
rect 15526 16838 15552 16890
rect 15256 16836 15312 16838
rect 15336 16836 15392 16838
rect 15416 16836 15472 16838
rect 15496 16836 15552 16838
rect 18256 16890 18312 16892
rect 18336 16890 18392 16892
rect 18416 16890 18472 16892
rect 18496 16890 18552 16892
rect 18256 16838 18282 16890
rect 18282 16838 18312 16890
rect 18336 16838 18346 16890
rect 18346 16838 18392 16890
rect 18416 16838 18462 16890
rect 18462 16838 18472 16890
rect 18496 16838 18526 16890
rect 18526 16838 18552 16890
rect 18256 16836 18312 16838
rect 18336 16836 18392 16838
rect 18416 16836 18472 16838
rect 18496 16836 18552 16838
rect 21256 16890 21312 16892
rect 21336 16890 21392 16892
rect 21416 16890 21472 16892
rect 21496 16890 21552 16892
rect 21256 16838 21282 16890
rect 21282 16838 21312 16890
rect 21336 16838 21346 16890
rect 21346 16838 21392 16890
rect 21416 16838 21462 16890
rect 21462 16838 21472 16890
rect 21496 16838 21526 16890
rect 21526 16838 21552 16890
rect 21256 16836 21312 16838
rect 21336 16836 21392 16838
rect 21416 16836 21472 16838
rect 21496 16836 21552 16838
rect 1756 16346 1812 16348
rect 1836 16346 1892 16348
rect 1916 16346 1972 16348
rect 1996 16346 2052 16348
rect 1756 16294 1782 16346
rect 1782 16294 1812 16346
rect 1836 16294 1846 16346
rect 1846 16294 1892 16346
rect 1916 16294 1962 16346
rect 1962 16294 1972 16346
rect 1996 16294 2026 16346
rect 2026 16294 2052 16346
rect 1756 16292 1812 16294
rect 1836 16292 1892 16294
rect 1916 16292 1972 16294
rect 1996 16292 2052 16294
rect 4756 16346 4812 16348
rect 4836 16346 4892 16348
rect 4916 16346 4972 16348
rect 4996 16346 5052 16348
rect 4756 16294 4782 16346
rect 4782 16294 4812 16346
rect 4836 16294 4846 16346
rect 4846 16294 4892 16346
rect 4916 16294 4962 16346
rect 4962 16294 4972 16346
rect 4996 16294 5026 16346
rect 5026 16294 5052 16346
rect 4756 16292 4812 16294
rect 4836 16292 4892 16294
rect 4916 16292 4972 16294
rect 4996 16292 5052 16294
rect 7756 16346 7812 16348
rect 7836 16346 7892 16348
rect 7916 16346 7972 16348
rect 7996 16346 8052 16348
rect 7756 16294 7782 16346
rect 7782 16294 7812 16346
rect 7836 16294 7846 16346
rect 7846 16294 7892 16346
rect 7916 16294 7962 16346
rect 7962 16294 7972 16346
rect 7996 16294 8026 16346
rect 8026 16294 8052 16346
rect 7756 16292 7812 16294
rect 7836 16292 7892 16294
rect 7916 16292 7972 16294
rect 7996 16292 8052 16294
rect 10756 16346 10812 16348
rect 10836 16346 10892 16348
rect 10916 16346 10972 16348
rect 10996 16346 11052 16348
rect 10756 16294 10782 16346
rect 10782 16294 10812 16346
rect 10836 16294 10846 16346
rect 10846 16294 10892 16346
rect 10916 16294 10962 16346
rect 10962 16294 10972 16346
rect 10996 16294 11026 16346
rect 11026 16294 11052 16346
rect 10756 16292 10812 16294
rect 10836 16292 10892 16294
rect 10916 16292 10972 16294
rect 10996 16292 11052 16294
rect 13756 16346 13812 16348
rect 13836 16346 13892 16348
rect 13916 16346 13972 16348
rect 13996 16346 14052 16348
rect 13756 16294 13782 16346
rect 13782 16294 13812 16346
rect 13836 16294 13846 16346
rect 13846 16294 13892 16346
rect 13916 16294 13962 16346
rect 13962 16294 13972 16346
rect 13996 16294 14026 16346
rect 14026 16294 14052 16346
rect 13756 16292 13812 16294
rect 13836 16292 13892 16294
rect 13916 16292 13972 16294
rect 13996 16292 14052 16294
rect 3256 15802 3312 15804
rect 3336 15802 3392 15804
rect 3416 15802 3472 15804
rect 3496 15802 3552 15804
rect 3256 15750 3282 15802
rect 3282 15750 3312 15802
rect 3336 15750 3346 15802
rect 3346 15750 3392 15802
rect 3416 15750 3462 15802
rect 3462 15750 3472 15802
rect 3496 15750 3526 15802
rect 3526 15750 3552 15802
rect 3256 15748 3312 15750
rect 3336 15748 3392 15750
rect 3416 15748 3472 15750
rect 3496 15748 3552 15750
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6416 15802 6472 15804
rect 6496 15802 6552 15804
rect 6256 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6416 15750 6462 15802
rect 6462 15750 6472 15802
rect 6496 15750 6526 15802
rect 6526 15750 6552 15802
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6416 15748 6472 15750
rect 6496 15748 6552 15750
rect 9256 15802 9312 15804
rect 9336 15802 9392 15804
rect 9416 15802 9472 15804
rect 9496 15802 9552 15804
rect 9256 15750 9282 15802
rect 9282 15750 9312 15802
rect 9336 15750 9346 15802
rect 9346 15750 9392 15802
rect 9416 15750 9462 15802
rect 9462 15750 9472 15802
rect 9496 15750 9526 15802
rect 9526 15750 9552 15802
rect 9256 15748 9312 15750
rect 9336 15748 9392 15750
rect 9416 15748 9472 15750
rect 9496 15748 9552 15750
rect 12256 15802 12312 15804
rect 12336 15802 12392 15804
rect 12416 15802 12472 15804
rect 12496 15802 12552 15804
rect 12256 15750 12282 15802
rect 12282 15750 12312 15802
rect 12336 15750 12346 15802
rect 12346 15750 12392 15802
rect 12416 15750 12462 15802
rect 12462 15750 12472 15802
rect 12496 15750 12526 15802
rect 12526 15750 12552 15802
rect 12256 15748 12312 15750
rect 12336 15748 12392 15750
rect 12416 15748 12472 15750
rect 12496 15748 12552 15750
rect 1756 15258 1812 15260
rect 1836 15258 1892 15260
rect 1916 15258 1972 15260
rect 1996 15258 2052 15260
rect 1756 15206 1782 15258
rect 1782 15206 1812 15258
rect 1836 15206 1846 15258
rect 1846 15206 1892 15258
rect 1916 15206 1962 15258
rect 1962 15206 1972 15258
rect 1996 15206 2026 15258
rect 2026 15206 2052 15258
rect 1756 15204 1812 15206
rect 1836 15204 1892 15206
rect 1916 15204 1972 15206
rect 1996 15204 2052 15206
rect 4756 15258 4812 15260
rect 4836 15258 4892 15260
rect 4916 15258 4972 15260
rect 4996 15258 5052 15260
rect 4756 15206 4782 15258
rect 4782 15206 4812 15258
rect 4836 15206 4846 15258
rect 4846 15206 4892 15258
rect 4916 15206 4962 15258
rect 4962 15206 4972 15258
rect 4996 15206 5026 15258
rect 5026 15206 5052 15258
rect 4756 15204 4812 15206
rect 4836 15204 4892 15206
rect 4916 15204 4972 15206
rect 4996 15204 5052 15206
rect 7756 15258 7812 15260
rect 7836 15258 7892 15260
rect 7916 15258 7972 15260
rect 7996 15258 8052 15260
rect 7756 15206 7782 15258
rect 7782 15206 7812 15258
rect 7836 15206 7846 15258
rect 7846 15206 7892 15258
rect 7916 15206 7962 15258
rect 7962 15206 7972 15258
rect 7996 15206 8026 15258
rect 8026 15206 8052 15258
rect 7756 15204 7812 15206
rect 7836 15204 7892 15206
rect 7916 15204 7972 15206
rect 7996 15204 8052 15206
rect 10756 15258 10812 15260
rect 10836 15258 10892 15260
rect 10916 15258 10972 15260
rect 10996 15258 11052 15260
rect 10756 15206 10782 15258
rect 10782 15206 10812 15258
rect 10836 15206 10846 15258
rect 10846 15206 10892 15258
rect 10916 15206 10962 15258
rect 10962 15206 10972 15258
rect 10996 15206 11026 15258
rect 11026 15206 11052 15258
rect 10756 15204 10812 15206
rect 10836 15204 10892 15206
rect 10916 15204 10972 15206
rect 10996 15204 11052 15206
rect 3256 14714 3312 14716
rect 3336 14714 3392 14716
rect 3416 14714 3472 14716
rect 3496 14714 3552 14716
rect 3256 14662 3282 14714
rect 3282 14662 3312 14714
rect 3336 14662 3346 14714
rect 3346 14662 3392 14714
rect 3416 14662 3462 14714
rect 3462 14662 3472 14714
rect 3496 14662 3526 14714
rect 3526 14662 3552 14714
rect 3256 14660 3312 14662
rect 3336 14660 3392 14662
rect 3416 14660 3472 14662
rect 3496 14660 3552 14662
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6416 14714 6472 14716
rect 6496 14714 6552 14716
rect 6256 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6416 14662 6462 14714
rect 6462 14662 6472 14714
rect 6496 14662 6526 14714
rect 6526 14662 6552 14714
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 6416 14660 6472 14662
rect 6496 14660 6552 14662
rect 9256 14714 9312 14716
rect 9336 14714 9392 14716
rect 9416 14714 9472 14716
rect 9496 14714 9552 14716
rect 9256 14662 9282 14714
rect 9282 14662 9312 14714
rect 9336 14662 9346 14714
rect 9346 14662 9392 14714
rect 9416 14662 9462 14714
rect 9462 14662 9472 14714
rect 9496 14662 9526 14714
rect 9526 14662 9552 14714
rect 9256 14660 9312 14662
rect 9336 14660 9392 14662
rect 9416 14660 9472 14662
rect 9496 14660 9552 14662
rect 12256 14714 12312 14716
rect 12336 14714 12392 14716
rect 12416 14714 12472 14716
rect 12496 14714 12552 14716
rect 12256 14662 12282 14714
rect 12282 14662 12312 14714
rect 12336 14662 12346 14714
rect 12346 14662 12392 14714
rect 12416 14662 12462 14714
rect 12462 14662 12472 14714
rect 12496 14662 12526 14714
rect 12526 14662 12552 14714
rect 12256 14660 12312 14662
rect 12336 14660 12392 14662
rect 12416 14660 12472 14662
rect 12496 14660 12552 14662
rect 1756 14170 1812 14172
rect 1836 14170 1892 14172
rect 1916 14170 1972 14172
rect 1996 14170 2052 14172
rect 1756 14118 1782 14170
rect 1782 14118 1812 14170
rect 1836 14118 1846 14170
rect 1846 14118 1892 14170
rect 1916 14118 1962 14170
rect 1962 14118 1972 14170
rect 1996 14118 2026 14170
rect 2026 14118 2052 14170
rect 1756 14116 1812 14118
rect 1836 14116 1892 14118
rect 1916 14116 1972 14118
rect 1996 14116 2052 14118
rect 4756 14170 4812 14172
rect 4836 14170 4892 14172
rect 4916 14170 4972 14172
rect 4996 14170 5052 14172
rect 4756 14118 4782 14170
rect 4782 14118 4812 14170
rect 4836 14118 4846 14170
rect 4846 14118 4892 14170
rect 4916 14118 4962 14170
rect 4962 14118 4972 14170
rect 4996 14118 5026 14170
rect 5026 14118 5052 14170
rect 4756 14116 4812 14118
rect 4836 14116 4892 14118
rect 4916 14116 4972 14118
rect 4996 14116 5052 14118
rect 7756 14170 7812 14172
rect 7836 14170 7892 14172
rect 7916 14170 7972 14172
rect 7996 14170 8052 14172
rect 7756 14118 7782 14170
rect 7782 14118 7812 14170
rect 7836 14118 7846 14170
rect 7846 14118 7892 14170
rect 7916 14118 7962 14170
rect 7962 14118 7972 14170
rect 7996 14118 8026 14170
rect 8026 14118 8052 14170
rect 7756 14116 7812 14118
rect 7836 14116 7892 14118
rect 7916 14116 7972 14118
rect 7996 14116 8052 14118
rect 10756 14170 10812 14172
rect 10836 14170 10892 14172
rect 10916 14170 10972 14172
rect 10996 14170 11052 14172
rect 10756 14118 10782 14170
rect 10782 14118 10812 14170
rect 10836 14118 10846 14170
rect 10846 14118 10892 14170
rect 10916 14118 10962 14170
rect 10962 14118 10972 14170
rect 10996 14118 11026 14170
rect 11026 14118 11052 14170
rect 10756 14116 10812 14118
rect 10836 14116 10892 14118
rect 10916 14116 10972 14118
rect 10996 14116 11052 14118
rect 13756 15258 13812 15260
rect 13836 15258 13892 15260
rect 13916 15258 13972 15260
rect 13996 15258 14052 15260
rect 13756 15206 13782 15258
rect 13782 15206 13812 15258
rect 13836 15206 13846 15258
rect 13846 15206 13892 15258
rect 13916 15206 13962 15258
rect 13962 15206 13972 15258
rect 13996 15206 14026 15258
rect 14026 15206 14052 15258
rect 13756 15204 13812 15206
rect 13836 15204 13892 15206
rect 13916 15204 13972 15206
rect 13996 15204 14052 15206
rect 15256 15802 15312 15804
rect 15336 15802 15392 15804
rect 15416 15802 15472 15804
rect 15496 15802 15552 15804
rect 15256 15750 15282 15802
rect 15282 15750 15312 15802
rect 15336 15750 15346 15802
rect 15346 15750 15392 15802
rect 15416 15750 15462 15802
rect 15462 15750 15472 15802
rect 15496 15750 15526 15802
rect 15526 15750 15552 15802
rect 15256 15748 15312 15750
rect 15336 15748 15392 15750
rect 15416 15748 15472 15750
rect 15496 15748 15552 15750
rect 110 13640 166 13696
rect 3256 13626 3312 13628
rect 3336 13626 3392 13628
rect 3416 13626 3472 13628
rect 3496 13626 3552 13628
rect 3256 13574 3282 13626
rect 3282 13574 3312 13626
rect 3336 13574 3346 13626
rect 3346 13574 3392 13626
rect 3416 13574 3462 13626
rect 3462 13574 3472 13626
rect 3496 13574 3526 13626
rect 3526 13574 3552 13626
rect 3256 13572 3312 13574
rect 3336 13572 3392 13574
rect 3416 13572 3472 13574
rect 3496 13572 3552 13574
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6416 13626 6472 13628
rect 6496 13626 6552 13628
rect 6256 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6416 13574 6462 13626
rect 6462 13574 6472 13626
rect 6496 13574 6526 13626
rect 6526 13574 6552 13626
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6416 13572 6472 13574
rect 6496 13572 6552 13574
rect 9256 13626 9312 13628
rect 9336 13626 9392 13628
rect 9416 13626 9472 13628
rect 9496 13626 9552 13628
rect 9256 13574 9282 13626
rect 9282 13574 9312 13626
rect 9336 13574 9346 13626
rect 9346 13574 9392 13626
rect 9416 13574 9462 13626
rect 9462 13574 9472 13626
rect 9496 13574 9526 13626
rect 9526 13574 9552 13626
rect 9256 13572 9312 13574
rect 9336 13572 9392 13574
rect 9416 13572 9472 13574
rect 9496 13572 9552 13574
rect 1756 13082 1812 13084
rect 1836 13082 1892 13084
rect 1916 13082 1972 13084
rect 1996 13082 2052 13084
rect 1756 13030 1782 13082
rect 1782 13030 1812 13082
rect 1836 13030 1846 13082
rect 1846 13030 1892 13082
rect 1916 13030 1962 13082
rect 1962 13030 1972 13082
rect 1996 13030 2026 13082
rect 2026 13030 2052 13082
rect 1756 13028 1812 13030
rect 1836 13028 1892 13030
rect 1916 13028 1972 13030
rect 1996 13028 2052 13030
rect 4756 13082 4812 13084
rect 4836 13082 4892 13084
rect 4916 13082 4972 13084
rect 4996 13082 5052 13084
rect 4756 13030 4782 13082
rect 4782 13030 4812 13082
rect 4836 13030 4846 13082
rect 4846 13030 4892 13082
rect 4916 13030 4962 13082
rect 4962 13030 4972 13082
rect 4996 13030 5026 13082
rect 5026 13030 5052 13082
rect 4756 13028 4812 13030
rect 4836 13028 4892 13030
rect 4916 13028 4972 13030
rect 4996 13028 5052 13030
rect 7756 13082 7812 13084
rect 7836 13082 7892 13084
rect 7916 13082 7972 13084
rect 7996 13082 8052 13084
rect 7756 13030 7782 13082
rect 7782 13030 7812 13082
rect 7836 13030 7846 13082
rect 7846 13030 7892 13082
rect 7916 13030 7962 13082
rect 7962 13030 7972 13082
rect 7996 13030 8026 13082
rect 8026 13030 8052 13082
rect 7756 13028 7812 13030
rect 7836 13028 7892 13030
rect 7916 13028 7972 13030
rect 7996 13028 8052 13030
rect 3256 12538 3312 12540
rect 3336 12538 3392 12540
rect 3416 12538 3472 12540
rect 3496 12538 3552 12540
rect 3256 12486 3282 12538
rect 3282 12486 3312 12538
rect 3336 12486 3346 12538
rect 3346 12486 3392 12538
rect 3416 12486 3462 12538
rect 3462 12486 3472 12538
rect 3496 12486 3526 12538
rect 3526 12486 3552 12538
rect 3256 12484 3312 12486
rect 3336 12484 3392 12486
rect 3416 12484 3472 12486
rect 3496 12484 3552 12486
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6416 12538 6472 12540
rect 6496 12538 6552 12540
rect 6256 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6416 12486 6462 12538
rect 6462 12486 6472 12538
rect 6496 12486 6526 12538
rect 6526 12486 6552 12538
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6416 12484 6472 12486
rect 6496 12484 6552 12486
rect 10756 13082 10812 13084
rect 10836 13082 10892 13084
rect 10916 13082 10972 13084
rect 10996 13082 11052 13084
rect 10756 13030 10782 13082
rect 10782 13030 10812 13082
rect 10836 13030 10846 13082
rect 10846 13030 10892 13082
rect 10916 13030 10962 13082
rect 10962 13030 10972 13082
rect 10996 13030 11026 13082
rect 11026 13030 11052 13082
rect 10756 13028 10812 13030
rect 10836 13028 10892 13030
rect 10916 13028 10972 13030
rect 10996 13028 11052 13030
rect 9256 12538 9312 12540
rect 9336 12538 9392 12540
rect 9416 12538 9472 12540
rect 9496 12538 9552 12540
rect 9256 12486 9282 12538
rect 9282 12486 9312 12538
rect 9336 12486 9346 12538
rect 9346 12486 9392 12538
rect 9416 12486 9462 12538
rect 9462 12486 9472 12538
rect 9496 12486 9526 12538
rect 9526 12486 9552 12538
rect 9256 12484 9312 12486
rect 9336 12484 9392 12486
rect 9416 12484 9472 12486
rect 9496 12484 9552 12486
rect 110 12144 166 12200
rect 1756 11994 1812 11996
rect 1836 11994 1892 11996
rect 1916 11994 1972 11996
rect 1996 11994 2052 11996
rect 1756 11942 1782 11994
rect 1782 11942 1812 11994
rect 1836 11942 1846 11994
rect 1846 11942 1892 11994
rect 1916 11942 1962 11994
rect 1962 11942 1972 11994
rect 1996 11942 2026 11994
rect 2026 11942 2052 11994
rect 1756 11940 1812 11942
rect 1836 11940 1892 11942
rect 1916 11940 1972 11942
rect 1996 11940 2052 11942
rect 4756 11994 4812 11996
rect 4836 11994 4892 11996
rect 4916 11994 4972 11996
rect 4996 11994 5052 11996
rect 4756 11942 4782 11994
rect 4782 11942 4812 11994
rect 4836 11942 4846 11994
rect 4846 11942 4892 11994
rect 4916 11942 4962 11994
rect 4962 11942 4972 11994
rect 4996 11942 5026 11994
rect 5026 11942 5052 11994
rect 4756 11940 4812 11942
rect 4836 11940 4892 11942
rect 4916 11940 4972 11942
rect 4996 11940 5052 11942
rect 7756 11994 7812 11996
rect 7836 11994 7892 11996
rect 7916 11994 7972 11996
rect 7996 11994 8052 11996
rect 7756 11942 7782 11994
rect 7782 11942 7812 11994
rect 7836 11942 7846 11994
rect 7846 11942 7892 11994
rect 7916 11942 7962 11994
rect 7962 11942 7972 11994
rect 7996 11942 8026 11994
rect 8026 11942 8052 11994
rect 7756 11940 7812 11942
rect 7836 11940 7892 11942
rect 7916 11940 7972 11942
rect 7996 11940 8052 11942
rect 3256 11450 3312 11452
rect 3336 11450 3392 11452
rect 3416 11450 3472 11452
rect 3496 11450 3552 11452
rect 3256 11398 3282 11450
rect 3282 11398 3312 11450
rect 3336 11398 3346 11450
rect 3346 11398 3392 11450
rect 3416 11398 3462 11450
rect 3462 11398 3472 11450
rect 3496 11398 3526 11450
rect 3526 11398 3552 11450
rect 3256 11396 3312 11398
rect 3336 11396 3392 11398
rect 3416 11396 3472 11398
rect 3496 11396 3552 11398
rect 1756 10906 1812 10908
rect 1836 10906 1892 10908
rect 1916 10906 1972 10908
rect 1996 10906 2052 10908
rect 1756 10854 1782 10906
rect 1782 10854 1812 10906
rect 1836 10854 1846 10906
rect 1846 10854 1892 10906
rect 1916 10854 1962 10906
rect 1962 10854 1972 10906
rect 1996 10854 2026 10906
rect 2026 10854 2052 10906
rect 1756 10852 1812 10854
rect 1836 10852 1892 10854
rect 1916 10852 1972 10854
rect 1996 10852 2052 10854
rect 4756 10906 4812 10908
rect 4836 10906 4892 10908
rect 4916 10906 4972 10908
rect 4996 10906 5052 10908
rect 4756 10854 4782 10906
rect 4782 10854 4812 10906
rect 4836 10854 4846 10906
rect 4846 10854 4892 10906
rect 4916 10854 4962 10906
rect 4962 10854 4972 10906
rect 4996 10854 5026 10906
rect 5026 10854 5052 10906
rect 4756 10852 4812 10854
rect 4836 10852 4892 10854
rect 4916 10852 4972 10854
rect 4996 10852 5052 10854
rect 3256 10362 3312 10364
rect 3336 10362 3392 10364
rect 3416 10362 3472 10364
rect 3496 10362 3552 10364
rect 3256 10310 3282 10362
rect 3282 10310 3312 10362
rect 3336 10310 3346 10362
rect 3346 10310 3392 10362
rect 3416 10310 3462 10362
rect 3462 10310 3472 10362
rect 3496 10310 3526 10362
rect 3526 10310 3552 10362
rect 3256 10308 3312 10310
rect 3336 10308 3392 10310
rect 3416 10308 3472 10310
rect 3496 10308 3552 10310
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6416 11450 6472 11452
rect 6496 11450 6552 11452
rect 6256 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6416 11398 6462 11450
rect 6462 11398 6472 11450
rect 6496 11398 6526 11450
rect 6526 11398 6552 11450
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6416 11396 6472 11398
rect 6496 11396 6552 11398
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6416 10362 6472 10364
rect 6496 10362 6552 10364
rect 6256 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6416 10310 6462 10362
rect 6462 10310 6472 10362
rect 6496 10310 6526 10362
rect 6526 10310 6552 10362
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6416 10308 6472 10310
rect 6496 10308 6552 10310
rect 7756 10906 7812 10908
rect 7836 10906 7892 10908
rect 7916 10906 7972 10908
rect 7996 10906 8052 10908
rect 7756 10854 7782 10906
rect 7782 10854 7812 10906
rect 7836 10854 7846 10906
rect 7846 10854 7892 10906
rect 7916 10854 7962 10906
rect 7962 10854 7972 10906
rect 7996 10854 8026 10906
rect 8026 10854 8052 10906
rect 7756 10852 7812 10854
rect 7836 10852 7892 10854
rect 7916 10852 7972 10854
rect 7996 10852 8052 10854
rect 1756 9818 1812 9820
rect 1836 9818 1892 9820
rect 1916 9818 1972 9820
rect 1996 9818 2052 9820
rect 1756 9766 1782 9818
rect 1782 9766 1812 9818
rect 1836 9766 1846 9818
rect 1846 9766 1892 9818
rect 1916 9766 1962 9818
rect 1962 9766 1972 9818
rect 1996 9766 2026 9818
rect 2026 9766 2052 9818
rect 1756 9764 1812 9766
rect 1836 9764 1892 9766
rect 1916 9764 1972 9766
rect 1996 9764 2052 9766
rect 4756 9818 4812 9820
rect 4836 9818 4892 9820
rect 4916 9818 4972 9820
rect 4996 9818 5052 9820
rect 4756 9766 4782 9818
rect 4782 9766 4812 9818
rect 4836 9766 4846 9818
rect 4846 9766 4892 9818
rect 4916 9766 4962 9818
rect 4962 9766 4972 9818
rect 4996 9766 5026 9818
rect 5026 9766 5052 9818
rect 4756 9764 4812 9766
rect 4836 9764 4892 9766
rect 4916 9764 4972 9766
rect 4996 9764 5052 9766
rect 3256 9274 3312 9276
rect 3336 9274 3392 9276
rect 3416 9274 3472 9276
rect 3496 9274 3552 9276
rect 3256 9222 3282 9274
rect 3282 9222 3312 9274
rect 3336 9222 3346 9274
rect 3346 9222 3392 9274
rect 3416 9222 3462 9274
rect 3462 9222 3472 9274
rect 3496 9222 3526 9274
rect 3526 9222 3552 9274
rect 3256 9220 3312 9222
rect 3336 9220 3392 9222
rect 3416 9220 3472 9222
rect 3496 9220 3552 9222
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6416 9274 6472 9276
rect 6496 9274 6552 9276
rect 6256 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6416 9222 6462 9274
rect 6462 9222 6472 9274
rect 6496 9222 6526 9274
rect 6526 9222 6552 9274
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 6416 9220 6472 9222
rect 6496 9220 6552 9222
rect 1756 8730 1812 8732
rect 1836 8730 1892 8732
rect 1916 8730 1972 8732
rect 1996 8730 2052 8732
rect 1756 8678 1782 8730
rect 1782 8678 1812 8730
rect 1836 8678 1846 8730
rect 1846 8678 1892 8730
rect 1916 8678 1962 8730
rect 1962 8678 1972 8730
rect 1996 8678 2026 8730
rect 2026 8678 2052 8730
rect 1756 8676 1812 8678
rect 1836 8676 1892 8678
rect 1916 8676 1972 8678
rect 1996 8676 2052 8678
rect 4756 8730 4812 8732
rect 4836 8730 4892 8732
rect 4916 8730 4972 8732
rect 4996 8730 5052 8732
rect 4756 8678 4782 8730
rect 4782 8678 4812 8730
rect 4836 8678 4846 8730
rect 4846 8678 4892 8730
rect 4916 8678 4962 8730
rect 4962 8678 4972 8730
rect 4996 8678 5026 8730
rect 5026 8678 5052 8730
rect 4756 8676 4812 8678
rect 4836 8676 4892 8678
rect 4916 8676 4972 8678
rect 4996 8676 5052 8678
rect 3256 8186 3312 8188
rect 3336 8186 3392 8188
rect 3416 8186 3472 8188
rect 3496 8186 3552 8188
rect 3256 8134 3282 8186
rect 3282 8134 3312 8186
rect 3336 8134 3346 8186
rect 3346 8134 3392 8186
rect 3416 8134 3462 8186
rect 3462 8134 3472 8186
rect 3496 8134 3526 8186
rect 3526 8134 3552 8186
rect 3256 8132 3312 8134
rect 3336 8132 3392 8134
rect 3416 8132 3472 8134
rect 3496 8132 3552 8134
rect 1756 7642 1812 7644
rect 1836 7642 1892 7644
rect 1916 7642 1972 7644
rect 1996 7642 2052 7644
rect 1756 7590 1782 7642
rect 1782 7590 1812 7642
rect 1836 7590 1846 7642
rect 1846 7590 1892 7642
rect 1916 7590 1962 7642
rect 1962 7590 1972 7642
rect 1996 7590 2026 7642
rect 2026 7590 2052 7642
rect 1756 7588 1812 7590
rect 1836 7588 1892 7590
rect 1916 7588 1972 7590
rect 1996 7588 2052 7590
rect 4756 7642 4812 7644
rect 4836 7642 4892 7644
rect 4916 7642 4972 7644
rect 4996 7642 5052 7644
rect 4756 7590 4782 7642
rect 4782 7590 4812 7642
rect 4836 7590 4846 7642
rect 4846 7590 4892 7642
rect 4916 7590 4962 7642
rect 4962 7590 4972 7642
rect 4996 7590 5026 7642
rect 5026 7590 5052 7642
rect 4756 7588 4812 7590
rect 4836 7588 4892 7590
rect 4916 7588 4972 7590
rect 4996 7588 5052 7590
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6416 8186 6472 8188
rect 6496 8186 6552 8188
rect 6256 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6416 8134 6462 8186
rect 6462 8134 6472 8186
rect 6496 8134 6526 8186
rect 6526 8134 6552 8186
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6416 8132 6472 8134
rect 6496 8132 6552 8134
rect 3256 7098 3312 7100
rect 3336 7098 3392 7100
rect 3416 7098 3472 7100
rect 3496 7098 3552 7100
rect 3256 7046 3282 7098
rect 3282 7046 3312 7098
rect 3336 7046 3346 7098
rect 3346 7046 3392 7098
rect 3416 7046 3462 7098
rect 3462 7046 3472 7098
rect 3496 7046 3526 7098
rect 3526 7046 3552 7098
rect 3256 7044 3312 7046
rect 3336 7044 3392 7046
rect 3416 7044 3472 7046
rect 3496 7044 3552 7046
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6416 7098 6472 7100
rect 6496 7098 6552 7100
rect 6256 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6416 7046 6462 7098
rect 6462 7046 6472 7098
rect 6496 7046 6526 7098
rect 6526 7046 6552 7098
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6416 7044 6472 7046
rect 6496 7044 6552 7046
rect 1756 6554 1812 6556
rect 1836 6554 1892 6556
rect 1916 6554 1972 6556
rect 1996 6554 2052 6556
rect 1756 6502 1782 6554
rect 1782 6502 1812 6554
rect 1836 6502 1846 6554
rect 1846 6502 1892 6554
rect 1916 6502 1962 6554
rect 1962 6502 1972 6554
rect 1996 6502 2026 6554
rect 2026 6502 2052 6554
rect 1756 6500 1812 6502
rect 1836 6500 1892 6502
rect 1916 6500 1972 6502
rect 1996 6500 2052 6502
rect 4756 6554 4812 6556
rect 4836 6554 4892 6556
rect 4916 6554 4972 6556
rect 4996 6554 5052 6556
rect 4756 6502 4782 6554
rect 4782 6502 4812 6554
rect 4836 6502 4846 6554
rect 4846 6502 4892 6554
rect 4916 6502 4962 6554
rect 4962 6502 4972 6554
rect 4996 6502 5026 6554
rect 5026 6502 5052 6554
rect 4756 6500 4812 6502
rect 4836 6500 4892 6502
rect 4916 6500 4972 6502
rect 4996 6500 5052 6502
rect 3256 6010 3312 6012
rect 3336 6010 3392 6012
rect 3416 6010 3472 6012
rect 3496 6010 3552 6012
rect 3256 5958 3282 6010
rect 3282 5958 3312 6010
rect 3336 5958 3346 6010
rect 3346 5958 3392 6010
rect 3416 5958 3462 6010
rect 3462 5958 3472 6010
rect 3496 5958 3526 6010
rect 3526 5958 3552 6010
rect 3256 5956 3312 5958
rect 3336 5956 3392 5958
rect 3416 5956 3472 5958
rect 3496 5956 3552 5958
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6416 6010 6472 6012
rect 6496 6010 6552 6012
rect 6256 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6416 5958 6462 6010
rect 6462 5958 6472 6010
rect 6496 5958 6526 6010
rect 6526 5958 6552 6010
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 6416 5956 6472 5958
rect 6496 5956 6552 5958
rect 7756 9818 7812 9820
rect 7836 9818 7892 9820
rect 7916 9818 7972 9820
rect 7996 9818 8052 9820
rect 7756 9766 7782 9818
rect 7782 9766 7812 9818
rect 7836 9766 7846 9818
rect 7846 9766 7892 9818
rect 7916 9766 7962 9818
rect 7962 9766 7972 9818
rect 7996 9766 8026 9818
rect 8026 9766 8052 9818
rect 7756 9764 7812 9766
rect 7836 9764 7892 9766
rect 7916 9764 7972 9766
rect 7996 9764 8052 9766
rect 7756 8730 7812 8732
rect 7836 8730 7892 8732
rect 7916 8730 7972 8732
rect 7996 8730 8052 8732
rect 7756 8678 7782 8730
rect 7782 8678 7812 8730
rect 7836 8678 7846 8730
rect 7846 8678 7892 8730
rect 7916 8678 7962 8730
rect 7962 8678 7972 8730
rect 7996 8678 8026 8730
rect 8026 8678 8052 8730
rect 7756 8676 7812 8678
rect 7836 8676 7892 8678
rect 7916 8676 7972 8678
rect 7996 8676 8052 8678
rect 7756 7642 7812 7644
rect 7836 7642 7892 7644
rect 7916 7642 7972 7644
rect 7996 7642 8052 7644
rect 7756 7590 7782 7642
rect 7782 7590 7812 7642
rect 7836 7590 7846 7642
rect 7846 7590 7892 7642
rect 7916 7590 7962 7642
rect 7962 7590 7972 7642
rect 7996 7590 8026 7642
rect 8026 7590 8052 7642
rect 7756 7588 7812 7590
rect 7836 7588 7892 7590
rect 7916 7588 7972 7590
rect 7996 7588 8052 7590
rect 7756 6554 7812 6556
rect 7836 6554 7892 6556
rect 7916 6554 7972 6556
rect 7996 6554 8052 6556
rect 7756 6502 7782 6554
rect 7782 6502 7812 6554
rect 7836 6502 7846 6554
rect 7846 6502 7892 6554
rect 7916 6502 7962 6554
rect 7962 6502 7972 6554
rect 7996 6502 8026 6554
rect 8026 6502 8052 6554
rect 7756 6500 7812 6502
rect 7836 6500 7892 6502
rect 7916 6500 7972 6502
rect 7996 6500 8052 6502
rect 10756 11994 10812 11996
rect 10836 11994 10892 11996
rect 10916 11994 10972 11996
rect 10996 11994 11052 11996
rect 10756 11942 10782 11994
rect 10782 11942 10812 11994
rect 10836 11942 10846 11994
rect 10846 11942 10892 11994
rect 10916 11942 10962 11994
rect 10962 11942 10972 11994
rect 10996 11942 11026 11994
rect 11026 11942 11052 11994
rect 10756 11940 10812 11942
rect 10836 11940 10892 11942
rect 10916 11940 10972 11942
rect 10996 11940 11052 11942
rect 9256 11450 9312 11452
rect 9336 11450 9392 11452
rect 9416 11450 9472 11452
rect 9496 11450 9552 11452
rect 9256 11398 9282 11450
rect 9282 11398 9312 11450
rect 9336 11398 9346 11450
rect 9346 11398 9392 11450
rect 9416 11398 9462 11450
rect 9462 11398 9472 11450
rect 9496 11398 9526 11450
rect 9526 11398 9552 11450
rect 9256 11396 9312 11398
rect 9336 11396 9392 11398
rect 9416 11396 9472 11398
rect 9496 11396 9552 11398
rect 9256 10362 9312 10364
rect 9336 10362 9392 10364
rect 9416 10362 9472 10364
rect 9496 10362 9552 10364
rect 9256 10310 9282 10362
rect 9282 10310 9312 10362
rect 9336 10310 9346 10362
rect 9346 10310 9392 10362
rect 9416 10310 9462 10362
rect 9462 10310 9472 10362
rect 9496 10310 9526 10362
rect 9526 10310 9552 10362
rect 9256 10308 9312 10310
rect 9336 10308 9392 10310
rect 9416 10308 9472 10310
rect 9496 10308 9552 10310
rect 12256 13626 12312 13628
rect 12336 13626 12392 13628
rect 12416 13626 12472 13628
rect 12496 13626 12552 13628
rect 12256 13574 12282 13626
rect 12282 13574 12312 13626
rect 12336 13574 12346 13626
rect 12346 13574 12392 13626
rect 12416 13574 12462 13626
rect 12462 13574 12472 13626
rect 12496 13574 12526 13626
rect 12526 13574 12552 13626
rect 12256 13572 12312 13574
rect 12336 13572 12392 13574
rect 12416 13572 12472 13574
rect 12496 13572 12552 13574
rect 13756 14170 13812 14172
rect 13836 14170 13892 14172
rect 13916 14170 13972 14172
rect 13996 14170 14052 14172
rect 13756 14118 13782 14170
rect 13782 14118 13812 14170
rect 13836 14118 13846 14170
rect 13846 14118 13892 14170
rect 13916 14118 13962 14170
rect 13962 14118 13972 14170
rect 13996 14118 14026 14170
rect 14026 14118 14052 14170
rect 13756 14116 13812 14118
rect 13836 14116 13892 14118
rect 13916 14116 13972 14118
rect 13996 14116 14052 14118
rect 15256 14714 15312 14716
rect 15336 14714 15392 14716
rect 15416 14714 15472 14716
rect 15496 14714 15552 14716
rect 15256 14662 15282 14714
rect 15282 14662 15312 14714
rect 15336 14662 15346 14714
rect 15346 14662 15392 14714
rect 15416 14662 15462 14714
rect 15462 14662 15472 14714
rect 15496 14662 15526 14714
rect 15526 14662 15552 14714
rect 15256 14660 15312 14662
rect 15336 14660 15392 14662
rect 15416 14660 15472 14662
rect 15496 14660 15552 14662
rect 12256 12538 12312 12540
rect 12336 12538 12392 12540
rect 12416 12538 12472 12540
rect 12496 12538 12552 12540
rect 12256 12486 12282 12538
rect 12282 12486 12312 12538
rect 12336 12486 12346 12538
rect 12346 12486 12392 12538
rect 12416 12486 12462 12538
rect 12462 12486 12472 12538
rect 12496 12486 12526 12538
rect 12526 12486 12552 12538
rect 12256 12484 12312 12486
rect 12336 12484 12392 12486
rect 12416 12484 12472 12486
rect 12496 12484 12552 12486
rect 10756 10906 10812 10908
rect 10836 10906 10892 10908
rect 10916 10906 10972 10908
rect 10996 10906 11052 10908
rect 10756 10854 10782 10906
rect 10782 10854 10812 10906
rect 10836 10854 10846 10906
rect 10846 10854 10892 10906
rect 10916 10854 10962 10906
rect 10962 10854 10972 10906
rect 10996 10854 11026 10906
rect 11026 10854 11052 10906
rect 10756 10852 10812 10854
rect 10836 10852 10892 10854
rect 10916 10852 10972 10854
rect 10996 10852 11052 10854
rect 9256 9274 9312 9276
rect 9336 9274 9392 9276
rect 9416 9274 9472 9276
rect 9496 9274 9552 9276
rect 9256 9222 9282 9274
rect 9282 9222 9312 9274
rect 9336 9222 9346 9274
rect 9346 9222 9392 9274
rect 9416 9222 9462 9274
rect 9462 9222 9472 9274
rect 9496 9222 9526 9274
rect 9526 9222 9552 9274
rect 9256 9220 9312 9222
rect 9336 9220 9392 9222
rect 9416 9220 9472 9222
rect 9496 9220 9552 9222
rect 9256 8186 9312 8188
rect 9336 8186 9392 8188
rect 9416 8186 9472 8188
rect 9496 8186 9552 8188
rect 9256 8134 9282 8186
rect 9282 8134 9312 8186
rect 9336 8134 9346 8186
rect 9346 8134 9392 8186
rect 9416 8134 9462 8186
rect 9462 8134 9472 8186
rect 9496 8134 9526 8186
rect 9526 8134 9552 8186
rect 9256 8132 9312 8134
rect 9336 8132 9392 8134
rect 9416 8132 9472 8134
rect 9496 8132 9552 8134
rect 9256 7098 9312 7100
rect 9336 7098 9392 7100
rect 9416 7098 9472 7100
rect 9496 7098 9552 7100
rect 9256 7046 9282 7098
rect 9282 7046 9312 7098
rect 9336 7046 9346 7098
rect 9346 7046 9392 7098
rect 9416 7046 9462 7098
rect 9462 7046 9472 7098
rect 9496 7046 9526 7098
rect 9526 7046 9552 7098
rect 9256 7044 9312 7046
rect 9336 7044 9392 7046
rect 9416 7044 9472 7046
rect 9496 7044 9552 7046
rect 10756 9818 10812 9820
rect 10836 9818 10892 9820
rect 10916 9818 10972 9820
rect 10996 9818 11052 9820
rect 10756 9766 10782 9818
rect 10782 9766 10812 9818
rect 10836 9766 10846 9818
rect 10846 9766 10892 9818
rect 10916 9766 10962 9818
rect 10962 9766 10972 9818
rect 10996 9766 11026 9818
rect 11026 9766 11052 9818
rect 10756 9764 10812 9766
rect 10836 9764 10892 9766
rect 10916 9764 10972 9766
rect 10996 9764 11052 9766
rect 12256 11450 12312 11452
rect 12336 11450 12392 11452
rect 12416 11450 12472 11452
rect 12496 11450 12552 11452
rect 12256 11398 12282 11450
rect 12282 11398 12312 11450
rect 12336 11398 12346 11450
rect 12346 11398 12392 11450
rect 12416 11398 12462 11450
rect 12462 11398 12472 11450
rect 12496 11398 12526 11450
rect 12526 11398 12552 11450
rect 12256 11396 12312 11398
rect 12336 11396 12392 11398
rect 12416 11396 12472 11398
rect 12496 11396 12552 11398
rect 13756 13082 13812 13084
rect 13836 13082 13892 13084
rect 13916 13082 13972 13084
rect 13996 13082 14052 13084
rect 13756 13030 13782 13082
rect 13782 13030 13812 13082
rect 13836 13030 13846 13082
rect 13846 13030 13892 13082
rect 13916 13030 13962 13082
rect 13962 13030 13972 13082
rect 13996 13030 14026 13082
rect 14026 13030 14052 13082
rect 13756 13028 13812 13030
rect 13836 13028 13892 13030
rect 13916 13028 13972 13030
rect 13996 13028 14052 13030
rect 13756 11994 13812 11996
rect 13836 11994 13892 11996
rect 13916 11994 13972 11996
rect 13996 11994 14052 11996
rect 13756 11942 13782 11994
rect 13782 11942 13812 11994
rect 13836 11942 13846 11994
rect 13846 11942 13892 11994
rect 13916 11942 13962 11994
rect 13962 11942 13972 11994
rect 13996 11942 14026 11994
rect 14026 11942 14052 11994
rect 13756 11940 13812 11942
rect 13836 11940 13892 11942
rect 13916 11940 13972 11942
rect 13996 11940 14052 11942
rect 15256 13626 15312 13628
rect 15336 13626 15392 13628
rect 15416 13626 15472 13628
rect 15496 13626 15552 13628
rect 15256 13574 15282 13626
rect 15282 13574 15312 13626
rect 15336 13574 15346 13626
rect 15346 13574 15392 13626
rect 15416 13574 15462 13626
rect 15462 13574 15472 13626
rect 15496 13574 15526 13626
rect 15526 13574 15552 13626
rect 15256 13572 15312 13574
rect 15336 13572 15392 13574
rect 15416 13572 15472 13574
rect 15496 13572 15552 13574
rect 12256 10362 12312 10364
rect 12336 10362 12392 10364
rect 12416 10362 12472 10364
rect 12496 10362 12552 10364
rect 12256 10310 12282 10362
rect 12282 10310 12312 10362
rect 12336 10310 12346 10362
rect 12346 10310 12392 10362
rect 12416 10310 12462 10362
rect 12462 10310 12472 10362
rect 12496 10310 12526 10362
rect 12526 10310 12552 10362
rect 12256 10308 12312 10310
rect 12336 10308 12392 10310
rect 12416 10308 12472 10310
rect 12496 10308 12552 10310
rect 10756 8730 10812 8732
rect 10836 8730 10892 8732
rect 10916 8730 10972 8732
rect 10996 8730 11052 8732
rect 10756 8678 10782 8730
rect 10782 8678 10812 8730
rect 10836 8678 10846 8730
rect 10846 8678 10892 8730
rect 10916 8678 10962 8730
rect 10962 8678 10972 8730
rect 10996 8678 11026 8730
rect 11026 8678 11052 8730
rect 10756 8676 10812 8678
rect 10836 8676 10892 8678
rect 10916 8676 10972 8678
rect 10996 8676 11052 8678
rect 10756 7642 10812 7644
rect 10836 7642 10892 7644
rect 10916 7642 10972 7644
rect 10996 7642 11052 7644
rect 10756 7590 10782 7642
rect 10782 7590 10812 7642
rect 10836 7590 10846 7642
rect 10846 7590 10892 7642
rect 10916 7590 10962 7642
rect 10962 7590 10972 7642
rect 10996 7590 11026 7642
rect 11026 7590 11052 7642
rect 10756 7588 10812 7590
rect 10836 7588 10892 7590
rect 10916 7588 10972 7590
rect 10996 7588 11052 7590
rect 1756 5466 1812 5468
rect 1836 5466 1892 5468
rect 1916 5466 1972 5468
rect 1996 5466 2052 5468
rect 1756 5414 1782 5466
rect 1782 5414 1812 5466
rect 1836 5414 1846 5466
rect 1846 5414 1892 5466
rect 1916 5414 1962 5466
rect 1962 5414 1972 5466
rect 1996 5414 2026 5466
rect 2026 5414 2052 5466
rect 1756 5412 1812 5414
rect 1836 5412 1892 5414
rect 1916 5412 1972 5414
rect 1996 5412 2052 5414
rect 4756 5466 4812 5468
rect 4836 5466 4892 5468
rect 4916 5466 4972 5468
rect 4996 5466 5052 5468
rect 4756 5414 4782 5466
rect 4782 5414 4812 5466
rect 4836 5414 4846 5466
rect 4846 5414 4892 5466
rect 4916 5414 4962 5466
rect 4962 5414 4972 5466
rect 4996 5414 5026 5466
rect 5026 5414 5052 5466
rect 4756 5412 4812 5414
rect 4836 5412 4892 5414
rect 4916 5412 4972 5414
rect 4996 5412 5052 5414
rect 3256 4922 3312 4924
rect 3336 4922 3392 4924
rect 3416 4922 3472 4924
rect 3496 4922 3552 4924
rect 3256 4870 3282 4922
rect 3282 4870 3312 4922
rect 3336 4870 3346 4922
rect 3346 4870 3392 4922
rect 3416 4870 3462 4922
rect 3462 4870 3472 4922
rect 3496 4870 3526 4922
rect 3526 4870 3552 4922
rect 3256 4868 3312 4870
rect 3336 4868 3392 4870
rect 3416 4868 3472 4870
rect 3496 4868 3552 4870
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6416 4922 6472 4924
rect 6496 4922 6552 4924
rect 6256 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6416 4870 6462 4922
rect 6462 4870 6472 4922
rect 6496 4870 6526 4922
rect 6526 4870 6552 4922
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 6416 4868 6472 4870
rect 6496 4868 6552 4870
rect 1756 4378 1812 4380
rect 1836 4378 1892 4380
rect 1916 4378 1972 4380
rect 1996 4378 2052 4380
rect 1756 4326 1782 4378
rect 1782 4326 1812 4378
rect 1836 4326 1846 4378
rect 1846 4326 1892 4378
rect 1916 4326 1962 4378
rect 1962 4326 1972 4378
rect 1996 4326 2026 4378
rect 2026 4326 2052 4378
rect 1756 4324 1812 4326
rect 1836 4324 1892 4326
rect 1916 4324 1972 4326
rect 1996 4324 2052 4326
rect 4756 4378 4812 4380
rect 4836 4378 4892 4380
rect 4916 4378 4972 4380
rect 4996 4378 5052 4380
rect 4756 4326 4782 4378
rect 4782 4326 4812 4378
rect 4836 4326 4846 4378
rect 4846 4326 4892 4378
rect 4916 4326 4962 4378
rect 4962 4326 4972 4378
rect 4996 4326 5026 4378
rect 5026 4326 5052 4378
rect 4756 4324 4812 4326
rect 4836 4324 4892 4326
rect 4916 4324 4972 4326
rect 4996 4324 5052 4326
rect 7756 5466 7812 5468
rect 7836 5466 7892 5468
rect 7916 5466 7972 5468
rect 7996 5466 8052 5468
rect 7756 5414 7782 5466
rect 7782 5414 7812 5466
rect 7836 5414 7846 5466
rect 7846 5414 7892 5466
rect 7916 5414 7962 5466
rect 7962 5414 7972 5466
rect 7996 5414 8026 5466
rect 8026 5414 8052 5466
rect 7756 5412 7812 5414
rect 7836 5412 7892 5414
rect 7916 5412 7972 5414
rect 7996 5412 8052 5414
rect 9256 6010 9312 6012
rect 9336 6010 9392 6012
rect 9416 6010 9472 6012
rect 9496 6010 9552 6012
rect 9256 5958 9282 6010
rect 9282 5958 9312 6010
rect 9336 5958 9346 6010
rect 9346 5958 9392 6010
rect 9416 5958 9462 6010
rect 9462 5958 9472 6010
rect 9496 5958 9526 6010
rect 9526 5958 9552 6010
rect 9256 5956 9312 5958
rect 9336 5956 9392 5958
rect 9416 5956 9472 5958
rect 9496 5956 9552 5958
rect 10756 6554 10812 6556
rect 10836 6554 10892 6556
rect 10916 6554 10972 6556
rect 10996 6554 11052 6556
rect 10756 6502 10782 6554
rect 10782 6502 10812 6554
rect 10836 6502 10846 6554
rect 10846 6502 10892 6554
rect 10916 6502 10962 6554
rect 10962 6502 10972 6554
rect 10996 6502 11026 6554
rect 11026 6502 11052 6554
rect 10756 6500 10812 6502
rect 10836 6500 10892 6502
rect 10916 6500 10972 6502
rect 10996 6500 11052 6502
rect 9256 4922 9312 4924
rect 9336 4922 9392 4924
rect 9416 4922 9472 4924
rect 9496 4922 9552 4924
rect 9256 4870 9282 4922
rect 9282 4870 9312 4922
rect 9336 4870 9346 4922
rect 9346 4870 9392 4922
rect 9416 4870 9462 4922
rect 9462 4870 9472 4922
rect 9496 4870 9526 4922
rect 9526 4870 9552 4922
rect 9256 4868 9312 4870
rect 9336 4868 9392 4870
rect 9416 4868 9472 4870
rect 9496 4868 9552 4870
rect 7756 4378 7812 4380
rect 7836 4378 7892 4380
rect 7916 4378 7972 4380
rect 7996 4378 8052 4380
rect 7756 4326 7782 4378
rect 7782 4326 7812 4378
rect 7836 4326 7846 4378
rect 7846 4326 7892 4378
rect 7916 4326 7962 4378
rect 7962 4326 7972 4378
rect 7996 4326 8026 4378
rect 8026 4326 8052 4378
rect 7756 4324 7812 4326
rect 7836 4324 7892 4326
rect 7916 4324 7972 4326
rect 7996 4324 8052 4326
rect 7654 3984 7710 4040
rect 3256 3834 3312 3836
rect 3336 3834 3392 3836
rect 3416 3834 3472 3836
rect 3496 3834 3552 3836
rect 3256 3782 3282 3834
rect 3282 3782 3312 3834
rect 3336 3782 3346 3834
rect 3346 3782 3392 3834
rect 3416 3782 3462 3834
rect 3462 3782 3472 3834
rect 3496 3782 3526 3834
rect 3526 3782 3552 3834
rect 3256 3780 3312 3782
rect 3336 3780 3392 3782
rect 3416 3780 3472 3782
rect 3496 3780 3552 3782
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6416 3834 6472 3836
rect 6496 3834 6552 3836
rect 6256 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6416 3782 6462 3834
rect 6462 3782 6472 3834
rect 6496 3782 6526 3834
rect 6526 3782 6552 3834
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 6416 3780 6472 3782
rect 6496 3780 6552 3782
rect 1756 3290 1812 3292
rect 1836 3290 1892 3292
rect 1916 3290 1972 3292
rect 1996 3290 2052 3292
rect 1756 3238 1782 3290
rect 1782 3238 1812 3290
rect 1836 3238 1846 3290
rect 1846 3238 1892 3290
rect 1916 3238 1962 3290
rect 1962 3238 1972 3290
rect 1996 3238 2026 3290
rect 2026 3238 2052 3290
rect 1756 3236 1812 3238
rect 1836 3236 1892 3238
rect 1916 3236 1972 3238
rect 1996 3236 2052 3238
rect 4756 3290 4812 3292
rect 4836 3290 4892 3292
rect 4916 3290 4972 3292
rect 4996 3290 5052 3292
rect 4756 3238 4782 3290
rect 4782 3238 4812 3290
rect 4836 3238 4846 3290
rect 4846 3238 4892 3290
rect 4916 3238 4962 3290
rect 4962 3238 4972 3290
rect 4996 3238 5026 3290
rect 5026 3238 5052 3290
rect 4756 3236 4812 3238
rect 4836 3236 4892 3238
rect 4916 3236 4972 3238
rect 4996 3236 5052 3238
rect 3256 2746 3312 2748
rect 3336 2746 3392 2748
rect 3416 2746 3472 2748
rect 3496 2746 3552 2748
rect 3256 2694 3282 2746
rect 3282 2694 3312 2746
rect 3336 2694 3346 2746
rect 3346 2694 3392 2746
rect 3416 2694 3462 2746
rect 3462 2694 3472 2746
rect 3496 2694 3526 2746
rect 3526 2694 3552 2746
rect 3256 2692 3312 2694
rect 3336 2692 3392 2694
rect 3416 2692 3472 2694
rect 3496 2692 3552 2694
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6416 2746 6472 2748
rect 6496 2746 6552 2748
rect 6256 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6416 2694 6462 2746
rect 6462 2694 6472 2746
rect 6496 2694 6526 2746
rect 6526 2694 6552 2746
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 6416 2692 6472 2694
rect 6496 2692 6552 2694
rect 7756 3290 7812 3292
rect 7836 3290 7892 3292
rect 7916 3290 7972 3292
rect 7996 3290 8052 3292
rect 7756 3238 7782 3290
rect 7782 3238 7812 3290
rect 7836 3238 7846 3290
rect 7846 3238 7892 3290
rect 7916 3238 7962 3290
rect 7962 3238 7972 3290
rect 7996 3238 8026 3290
rect 8026 3238 8052 3290
rect 7756 3236 7812 3238
rect 7836 3236 7892 3238
rect 7916 3236 7972 3238
rect 7996 3236 8052 3238
rect 9256 3834 9312 3836
rect 9336 3834 9392 3836
rect 9416 3834 9472 3836
rect 9496 3834 9552 3836
rect 9256 3782 9282 3834
rect 9282 3782 9312 3834
rect 9336 3782 9346 3834
rect 9346 3782 9392 3834
rect 9416 3782 9462 3834
rect 9462 3782 9472 3834
rect 9496 3782 9526 3834
rect 9526 3782 9552 3834
rect 9256 3780 9312 3782
rect 9336 3780 9392 3782
rect 9416 3780 9472 3782
rect 9496 3780 9552 3782
rect 9256 2746 9312 2748
rect 9336 2746 9392 2748
rect 9416 2746 9472 2748
rect 9496 2746 9552 2748
rect 9256 2694 9282 2746
rect 9282 2694 9312 2746
rect 9336 2694 9346 2746
rect 9346 2694 9392 2746
rect 9416 2694 9462 2746
rect 9462 2694 9472 2746
rect 9496 2694 9526 2746
rect 9526 2694 9552 2746
rect 9256 2692 9312 2694
rect 9336 2692 9392 2694
rect 9416 2692 9472 2694
rect 9496 2692 9552 2694
rect 1756 2202 1812 2204
rect 1836 2202 1892 2204
rect 1916 2202 1972 2204
rect 1996 2202 2052 2204
rect 1756 2150 1782 2202
rect 1782 2150 1812 2202
rect 1836 2150 1846 2202
rect 1846 2150 1892 2202
rect 1916 2150 1962 2202
rect 1962 2150 1972 2202
rect 1996 2150 2026 2202
rect 2026 2150 2052 2202
rect 1756 2148 1812 2150
rect 1836 2148 1892 2150
rect 1916 2148 1972 2150
rect 1996 2148 2052 2150
rect 4756 2202 4812 2204
rect 4836 2202 4892 2204
rect 4916 2202 4972 2204
rect 4996 2202 5052 2204
rect 4756 2150 4782 2202
rect 4782 2150 4812 2202
rect 4836 2150 4846 2202
rect 4846 2150 4892 2202
rect 4916 2150 4962 2202
rect 4962 2150 4972 2202
rect 4996 2150 5026 2202
rect 5026 2150 5052 2202
rect 4756 2148 4812 2150
rect 4836 2148 4892 2150
rect 4916 2148 4972 2150
rect 4996 2148 5052 2150
rect 7756 2202 7812 2204
rect 7836 2202 7892 2204
rect 7916 2202 7972 2204
rect 7996 2202 8052 2204
rect 7756 2150 7782 2202
rect 7782 2150 7812 2202
rect 7836 2150 7846 2202
rect 7846 2150 7892 2202
rect 7916 2150 7962 2202
rect 7962 2150 7972 2202
rect 7996 2150 8026 2202
rect 8026 2150 8052 2202
rect 7756 2148 7812 2150
rect 7836 2148 7892 2150
rect 7916 2148 7972 2150
rect 7996 2148 8052 2150
rect 10756 5466 10812 5468
rect 10836 5466 10892 5468
rect 10916 5466 10972 5468
rect 10996 5466 11052 5468
rect 10756 5414 10782 5466
rect 10782 5414 10812 5466
rect 10836 5414 10846 5466
rect 10846 5414 10892 5466
rect 10916 5414 10962 5466
rect 10962 5414 10972 5466
rect 10996 5414 11026 5466
rect 11026 5414 11052 5466
rect 10756 5412 10812 5414
rect 10836 5412 10892 5414
rect 10916 5412 10972 5414
rect 10996 5412 11052 5414
rect 13756 10906 13812 10908
rect 13836 10906 13892 10908
rect 13916 10906 13972 10908
rect 13996 10906 14052 10908
rect 13756 10854 13782 10906
rect 13782 10854 13812 10906
rect 13836 10854 13846 10906
rect 13846 10854 13892 10906
rect 13916 10854 13962 10906
rect 13962 10854 13972 10906
rect 13996 10854 14026 10906
rect 14026 10854 14052 10906
rect 13756 10852 13812 10854
rect 13836 10852 13892 10854
rect 13916 10852 13972 10854
rect 13996 10852 14052 10854
rect 13756 9818 13812 9820
rect 13836 9818 13892 9820
rect 13916 9818 13972 9820
rect 13996 9818 14052 9820
rect 13756 9766 13782 9818
rect 13782 9766 13812 9818
rect 13836 9766 13846 9818
rect 13846 9766 13892 9818
rect 13916 9766 13962 9818
rect 13962 9766 13972 9818
rect 13996 9766 14026 9818
rect 14026 9766 14052 9818
rect 13756 9764 13812 9766
rect 13836 9764 13892 9766
rect 13916 9764 13972 9766
rect 13996 9764 14052 9766
rect 12256 9274 12312 9276
rect 12336 9274 12392 9276
rect 12416 9274 12472 9276
rect 12496 9274 12552 9276
rect 12256 9222 12282 9274
rect 12282 9222 12312 9274
rect 12336 9222 12346 9274
rect 12346 9222 12392 9274
rect 12416 9222 12462 9274
rect 12462 9222 12472 9274
rect 12496 9222 12526 9274
rect 12526 9222 12552 9274
rect 12256 9220 12312 9222
rect 12336 9220 12392 9222
rect 12416 9220 12472 9222
rect 12496 9220 12552 9222
rect 12256 8186 12312 8188
rect 12336 8186 12392 8188
rect 12416 8186 12472 8188
rect 12496 8186 12552 8188
rect 12256 8134 12282 8186
rect 12282 8134 12312 8186
rect 12336 8134 12346 8186
rect 12346 8134 12392 8186
rect 12416 8134 12462 8186
rect 12462 8134 12472 8186
rect 12496 8134 12526 8186
rect 12526 8134 12552 8186
rect 12256 8132 12312 8134
rect 12336 8132 12392 8134
rect 12416 8132 12472 8134
rect 12496 8132 12552 8134
rect 10756 4378 10812 4380
rect 10836 4378 10892 4380
rect 10916 4378 10972 4380
rect 10996 4378 11052 4380
rect 10756 4326 10782 4378
rect 10782 4326 10812 4378
rect 10836 4326 10846 4378
rect 10846 4326 10892 4378
rect 10916 4326 10962 4378
rect 10962 4326 10972 4378
rect 10996 4326 11026 4378
rect 11026 4326 11052 4378
rect 10756 4324 10812 4326
rect 10836 4324 10892 4326
rect 10916 4324 10972 4326
rect 10996 4324 11052 4326
rect 10046 3984 10102 4040
rect 10756 3290 10812 3292
rect 10836 3290 10892 3292
rect 10916 3290 10972 3292
rect 10996 3290 11052 3292
rect 10756 3238 10782 3290
rect 10782 3238 10812 3290
rect 10836 3238 10846 3290
rect 10846 3238 10892 3290
rect 10916 3238 10962 3290
rect 10962 3238 10972 3290
rect 10996 3238 11026 3290
rect 11026 3238 11052 3290
rect 10756 3236 10812 3238
rect 10836 3236 10892 3238
rect 10916 3236 10972 3238
rect 10996 3236 11052 3238
rect 10046 2488 10102 2544
rect 12256 7098 12312 7100
rect 12336 7098 12392 7100
rect 12416 7098 12472 7100
rect 12496 7098 12552 7100
rect 12256 7046 12282 7098
rect 12282 7046 12312 7098
rect 12336 7046 12346 7098
rect 12346 7046 12392 7098
rect 12416 7046 12462 7098
rect 12462 7046 12472 7098
rect 12496 7046 12526 7098
rect 12526 7046 12552 7098
rect 12256 7044 12312 7046
rect 12336 7044 12392 7046
rect 12416 7044 12472 7046
rect 12496 7044 12552 7046
rect 13756 8730 13812 8732
rect 13836 8730 13892 8732
rect 13916 8730 13972 8732
rect 13996 8730 14052 8732
rect 13756 8678 13782 8730
rect 13782 8678 13812 8730
rect 13836 8678 13846 8730
rect 13846 8678 13892 8730
rect 13916 8678 13962 8730
rect 13962 8678 13972 8730
rect 13996 8678 14026 8730
rect 14026 8678 14052 8730
rect 13756 8676 13812 8678
rect 13836 8676 13892 8678
rect 13916 8676 13972 8678
rect 13996 8676 14052 8678
rect 13756 7642 13812 7644
rect 13836 7642 13892 7644
rect 13916 7642 13972 7644
rect 13996 7642 14052 7644
rect 13756 7590 13782 7642
rect 13782 7590 13812 7642
rect 13836 7590 13846 7642
rect 13846 7590 13892 7642
rect 13916 7590 13962 7642
rect 13962 7590 13972 7642
rect 13996 7590 14026 7642
rect 14026 7590 14052 7642
rect 13756 7588 13812 7590
rect 13836 7588 13892 7590
rect 13916 7588 13972 7590
rect 13996 7588 14052 7590
rect 13756 6554 13812 6556
rect 13836 6554 13892 6556
rect 13916 6554 13972 6556
rect 13996 6554 14052 6556
rect 13756 6502 13782 6554
rect 13782 6502 13812 6554
rect 13836 6502 13846 6554
rect 13846 6502 13892 6554
rect 13916 6502 13962 6554
rect 13962 6502 13972 6554
rect 13996 6502 14026 6554
rect 14026 6502 14052 6554
rect 13756 6500 13812 6502
rect 13836 6500 13892 6502
rect 13916 6500 13972 6502
rect 13996 6500 14052 6502
rect 12256 6010 12312 6012
rect 12336 6010 12392 6012
rect 12416 6010 12472 6012
rect 12496 6010 12552 6012
rect 12256 5958 12282 6010
rect 12282 5958 12312 6010
rect 12336 5958 12346 6010
rect 12346 5958 12392 6010
rect 12416 5958 12462 6010
rect 12462 5958 12472 6010
rect 12496 5958 12526 6010
rect 12526 5958 12552 6010
rect 12256 5956 12312 5958
rect 12336 5956 12392 5958
rect 12416 5956 12472 5958
rect 12496 5956 12552 5958
rect 12256 4922 12312 4924
rect 12336 4922 12392 4924
rect 12416 4922 12472 4924
rect 12496 4922 12552 4924
rect 12256 4870 12282 4922
rect 12282 4870 12312 4922
rect 12336 4870 12346 4922
rect 12346 4870 12392 4922
rect 12416 4870 12462 4922
rect 12462 4870 12472 4922
rect 12496 4870 12526 4922
rect 12526 4870 12552 4922
rect 12256 4868 12312 4870
rect 12336 4868 12392 4870
rect 12416 4868 12472 4870
rect 12496 4868 12552 4870
rect 12256 3834 12312 3836
rect 12336 3834 12392 3836
rect 12416 3834 12472 3836
rect 12496 3834 12552 3836
rect 12256 3782 12282 3834
rect 12282 3782 12312 3834
rect 12336 3782 12346 3834
rect 12346 3782 12392 3834
rect 12416 3782 12462 3834
rect 12462 3782 12472 3834
rect 12496 3782 12526 3834
rect 12526 3782 12552 3834
rect 12256 3780 12312 3782
rect 12336 3780 12392 3782
rect 12416 3780 12472 3782
rect 12496 3780 12552 3782
rect 12256 2746 12312 2748
rect 12336 2746 12392 2748
rect 12416 2746 12472 2748
rect 12496 2746 12552 2748
rect 12256 2694 12282 2746
rect 12282 2694 12312 2746
rect 12336 2694 12346 2746
rect 12346 2694 12392 2746
rect 12416 2694 12462 2746
rect 12462 2694 12472 2746
rect 12496 2694 12526 2746
rect 12526 2694 12552 2746
rect 12256 2692 12312 2694
rect 12336 2692 12392 2694
rect 12416 2692 12472 2694
rect 12496 2692 12552 2694
rect 13756 5466 13812 5468
rect 13836 5466 13892 5468
rect 13916 5466 13972 5468
rect 13996 5466 14052 5468
rect 13756 5414 13782 5466
rect 13782 5414 13812 5466
rect 13836 5414 13846 5466
rect 13846 5414 13892 5466
rect 13916 5414 13962 5466
rect 13962 5414 13972 5466
rect 13996 5414 14026 5466
rect 14026 5414 14052 5466
rect 13756 5412 13812 5414
rect 13836 5412 13892 5414
rect 13916 5412 13972 5414
rect 13996 5412 14052 5414
rect 15256 12538 15312 12540
rect 15336 12538 15392 12540
rect 15416 12538 15472 12540
rect 15496 12538 15552 12540
rect 15256 12486 15282 12538
rect 15282 12486 15312 12538
rect 15336 12486 15346 12538
rect 15346 12486 15392 12538
rect 15416 12486 15462 12538
rect 15462 12486 15472 12538
rect 15496 12486 15526 12538
rect 15526 12486 15552 12538
rect 15256 12484 15312 12486
rect 15336 12484 15392 12486
rect 15416 12484 15472 12486
rect 15496 12484 15552 12486
rect 15256 11450 15312 11452
rect 15336 11450 15392 11452
rect 15416 11450 15472 11452
rect 15496 11450 15552 11452
rect 15256 11398 15282 11450
rect 15282 11398 15312 11450
rect 15336 11398 15346 11450
rect 15346 11398 15392 11450
rect 15416 11398 15462 11450
rect 15462 11398 15472 11450
rect 15496 11398 15526 11450
rect 15526 11398 15552 11450
rect 15256 11396 15312 11398
rect 15336 11396 15392 11398
rect 15416 11396 15472 11398
rect 15496 11396 15552 11398
rect 16756 16346 16812 16348
rect 16836 16346 16892 16348
rect 16916 16346 16972 16348
rect 16996 16346 17052 16348
rect 16756 16294 16782 16346
rect 16782 16294 16812 16346
rect 16836 16294 16846 16346
rect 16846 16294 16892 16346
rect 16916 16294 16962 16346
rect 16962 16294 16972 16346
rect 16996 16294 17026 16346
rect 17026 16294 17052 16346
rect 16756 16292 16812 16294
rect 16836 16292 16892 16294
rect 16916 16292 16972 16294
rect 16996 16292 17052 16294
rect 19756 16346 19812 16348
rect 19836 16346 19892 16348
rect 19916 16346 19972 16348
rect 19996 16346 20052 16348
rect 19756 16294 19782 16346
rect 19782 16294 19812 16346
rect 19836 16294 19846 16346
rect 19846 16294 19892 16346
rect 19916 16294 19962 16346
rect 19962 16294 19972 16346
rect 19996 16294 20026 16346
rect 20026 16294 20052 16346
rect 19756 16292 19812 16294
rect 19836 16292 19892 16294
rect 19916 16292 19972 16294
rect 19996 16292 20052 16294
rect 18256 15802 18312 15804
rect 18336 15802 18392 15804
rect 18416 15802 18472 15804
rect 18496 15802 18552 15804
rect 18256 15750 18282 15802
rect 18282 15750 18312 15802
rect 18336 15750 18346 15802
rect 18346 15750 18392 15802
rect 18416 15750 18462 15802
rect 18462 15750 18472 15802
rect 18496 15750 18526 15802
rect 18526 15750 18552 15802
rect 18256 15748 18312 15750
rect 18336 15748 18392 15750
rect 18416 15748 18472 15750
rect 18496 15748 18552 15750
rect 21256 15802 21312 15804
rect 21336 15802 21392 15804
rect 21416 15802 21472 15804
rect 21496 15802 21552 15804
rect 21256 15750 21282 15802
rect 21282 15750 21312 15802
rect 21336 15750 21346 15802
rect 21346 15750 21392 15802
rect 21416 15750 21462 15802
rect 21462 15750 21472 15802
rect 21496 15750 21526 15802
rect 21526 15750 21552 15802
rect 21256 15748 21312 15750
rect 21336 15748 21392 15750
rect 21416 15748 21472 15750
rect 21496 15748 21552 15750
rect 16756 15258 16812 15260
rect 16836 15258 16892 15260
rect 16916 15258 16972 15260
rect 16996 15258 17052 15260
rect 16756 15206 16782 15258
rect 16782 15206 16812 15258
rect 16836 15206 16846 15258
rect 16846 15206 16892 15258
rect 16916 15206 16962 15258
rect 16962 15206 16972 15258
rect 16996 15206 17026 15258
rect 17026 15206 17052 15258
rect 16756 15204 16812 15206
rect 16836 15204 16892 15206
rect 16916 15204 16972 15206
rect 16996 15204 17052 15206
rect 16756 14170 16812 14172
rect 16836 14170 16892 14172
rect 16916 14170 16972 14172
rect 16996 14170 17052 14172
rect 16756 14118 16782 14170
rect 16782 14118 16812 14170
rect 16836 14118 16846 14170
rect 16846 14118 16892 14170
rect 16916 14118 16962 14170
rect 16962 14118 16972 14170
rect 16996 14118 17026 14170
rect 17026 14118 17052 14170
rect 16756 14116 16812 14118
rect 16836 14116 16892 14118
rect 16916 14116 16972 14118
rect 16996 14116 17052 14118
rect 18256 14714 18312 14716
rect 18336 14714 18392 14716
rect 18416 14714 18472 14716
rect 18496 14714 18552 14716
rect 18256 14662 18282 14714
rect 18282 14662 18312 14714
rect 18336 14662 18346 14714
rect 18346 14662 18392 14714
rect 18416 14662 18462 14714
rect 18462 14662 18472 14714
rect 18496 14662 18526 14714
rect 18526 14662 18552 14714
rect 18256 14660 18312 14662
rect 18336 14660 18392 14662
rect 18416 14660 18472 14662
rect 18496 14660 18552 14662
rect 16756 13082 16812 13084
rect 16836 13082 16892 13084
rect 16916 13082 16972 13084
rect 16996 13082 17052 13084
rect 16756 13030 16782 13082
rect 16782 13030 16812 13082
rect 16836 13030 16846 13082
rect 16846 13030 16892 13082
rect 16916 13030 16962 13082
rect 16962 13030 16972 13082
rect 16996 13030 17026 13082
rect 17026 13030 17052 13082
rect 16756 13028 16812 13030
rect 16836 13028 16892 13030
rect 16916 13028 16972 13030
rect 16996 13028 17052 13030
rect 18256 13626 18312 13628
rect 18336 13626 18392 13628
rect 18416 13626 18472 13628
rect 18496 13626 18552 13628
rect 18256 13574 18282 13626
rect 18282 13574 18312 13626
rect 18336 13574 18346 13626
rect 18346 13574 18392 13626
rect 18416 13574 18462 13626
rect 18462 13574 18472 13626
rect 18496 13574 18526 13626
rect 18526 13574 18552 13626
rect 18256 13572 18312 13574
rect 18336 13572 18392 13574
rect 18416 13572 18472 13574
rect 18496 13572 18552 13574
rect 19756 15258 19812 15260
rect 19836 15258 19892 15260
rect 19916 15258 19972 15260
rect 19996 15258 20052 15260
rect 19756 15206 19782 15258
rect 19782 15206 19812 15258
rect 19836 15206 19846 15258
rect 19846 15206 19892 15258
rect 19916 15206 19962 15258
rect 19962 15206 19972 15258
rect 19996 15206 20026 15258
rect 20026 15206 20052 15258
rect 19756 15204 19812 15206
rect 19836 15204 19892 15206
rect 19916 15204 19972 15206
rect 19996 15204 20052 15206
rect 19756 14170 19812 14172
rect 19836 14170 19892 14172
rect 19916 14170 19972 14172
rect 19996 14170 20052 14172
rect 19756 14118 19782 14170
rect 19782 14118 19812 14170
rect 19836 14118 19846 14170
rect 19846 14118 19892 14170
rect 19916 14118 19962 14170
rect 19962 14118 19972 14170
rect 19996 14118 20026 14170
rect 20026 14118 20052 14170
rect 19756 14116 19812 14118
rect 19836 14116 19892 14118
rect 19916 14116 19972 14118
rect 19996 14116 20052 14118
rect 15256 10362 15312 10364
rect 15336 10362 15392 10364
rect 15416 10362 15472 10364
rect 15496 10362 15552 10364
rect 15256 10310 15282 10362
rect 15282 10310 15312 10362
rect 15336 10310 15346 10362
rect 15346 10310 15392 10362
rect 15416 10310 15462 10362
rect 15462 10310 15472 10362
rect 15496 10310 15526 10362
rect 15526 10310 15552 10362
rect 15256 10308 15312 10310
rect 15336 10308 15392 10310
rect 15416 10308 15472 10310
rect 15496 10308 15552 10310
rect 15256 9274 15312 9276
rect 15336 9274 15392 9276
rect 15416 9274 15472 9276
rect 15496 9274 15552 9276
rect 15256 9222 15282 9274
rect 15282 9222 15312 9274
rect 15336 9222 15346 9274
rect 15346 9222 15392 9274
rect 15416 9222 15462 9274
rect 15462 9222 15472 9274
rect 15496 9222 15526 9274
rect 15526 9222 15552 9274
rect 15256 9220 15312 9222
rect 15336 9220 15392 9222
rect 15416 9220 15472 9222
rect 15496 9220 15552 9222
rect 15256 8186 15312 8188
rect 15336 8186 15392 8188
rect 15416 8186 15472 8188
rect 15496 8186 15552 8188
rect 15256 8134 15282 8186
rect 15282 8134 15312 8186
rect 15336 8134 15346 8186
rect 15346 8134 15392 8186
rect 15416 8134 15462 8186
rect 15462 8134 15472 8186
rect 15496 8134 15526 8186
rect 15526 8134 15552 8186
rect 15256 8132 15312 8134
rect 15336 8132 15392 8134
rect 15416 8132 15472 8134
rect 15496 8132 15552 8134
rect 15256 7098 15312 7100
rect 15336 7098 15392 7100
rect 15416 7098 15472 7100
rect 15496 7098 15552 7100
rect 15256 7046 15282 7098
rect 15282 7046 15312 7098
rect 15336 7046 15346 7098
rect 15346 7046 15392 7098
rect 15416 7046 15462 7098
rect 15462 7046 15472 7098
rect 15496 7046 15526 7098
rect 15526 7046 15552 7098
rect 15256 7044 15312 7046
rect 15336 7044 15392 7046
rect 15416 7044 15472 7046
rect 15496 7044 15552 7046
rect 16756 11994 16812 11996
rect 16836 11994 16892 11996
rect 16916 11994 16972 11996
rect 16996 11994 17052 11996
rect 16756 11942 16782 11994
rect 16782 11942 16812 11994
rect 16836 11942 16846 11994
rect 16846 11942 16892 11994
rect 16916 11942 16962 11994
rect 16962 11942 16972 11994
rect 16996 11942 17026 11994
rect 17026 11942 17052 11994
rect 16756 11940 16812 11942
rect 16836 11940 16892 11942
rect 16916 11940 16972 11942
rect 16996 11940 17052 11942
rect 16756 10906 16812 10908
rect 16836 10906 16892 10908
rect 16916 10906 16972 10908
rect 16996 10906 17052 10908
rect 16756 10854 16782 10906
rect 16782 10854 16812 10906
rect 16836 10854 16846 10906
rect 16846 10854 16892 10906
rect 16916 10854 16962 10906
rect 16962 10854 16972 10906
rect 16996 10854 17026 10906
rect 17026 10854 17052 10906
rect 16756 10852 16812 10854
rect 16836 10852 16892 10854
rect 16916 10852 16972 10854
rect 16996 10852 17052 10854
rect 16756 9818 16812 9820
rect 16836 9818 16892 9820
rect 16916 9818 16972 9820
rect 16996 9818 17052 9820
rect 16756 9766 16782 9818
rect 16782 9766 16812 9818
rect 16836 9766 16846 9818
rect 16846 9766 16892 9818
rect 16916 9766 16962 9818
rect 16962 9766 16972 9818
rect 16996 9766 17026 9818
rect 17026 9766 17052 9818
rect 16756 9764 16812 9766
rect 16836 9764 16892 9766
rect 16916 9764 16972 9766
rect 16996 9764 17052 9766
rect 18256 12538 18312 12540
rect 18336 12538 18392 12540
rect 18416 12538 18472 12540
rect 18496 12538 18552 12540
rect 18256 12486 18282 12538
rect 18282 12486 18312 12538
rect 18336 12486 18346 12538
rect 18346 12486 18392 12538
rect 18416 12486 18462 12538
rect 18462 12486 18472 12538
rect 18496 12486 18526 12538
rect 18526 12486 18552 12538
rect 18256 12484 18312 12486
rect 18336 12484 18392 12486
rect 18416 12484 18472 12486
rect 18496 12484 18552 12486
rect 18418 11736 18474 11792
rect 18256 11450 18312 11452
rect 18336 11450 18392 11452
rect 18416 11450 18472 11452
rect 18496 11450 18552 11452
rect 18256 11398 18282 11450
rect 18282 11398 18312 11450
rect 18336 11398 18346 11450
rect 18346 11398 18392 11450
rect 18416 11398 18462 11450
rect 18462 11398 18472 11450
rect 18496 11398 18526 11450
rect 18526 11398 18552 11450
rect 18256 11396 18312 11398
rect 18336 11396 18392 11398
rect 18416 11396 18472 11398
rect 18496 11396 18552 11398
rect 18256 10362 18312 10364
rect 18336 10362 18392 10364
rect 18416 10362 18472 10364
rect 18496 10362 18552 10364
rect 18256 10310 18282 10362
rect 18282 10310 18312 10362
rect 18336 10310 18346 10362
rect 18346 10310 18392 10362
rect 18416 10310 18462 10362
rect 18462 10310 18472 10362
rect 18496 10310 18526 10362
rect 18526 10310 18552 10362
rect 18256 10308 18312 10310
rect 18336 10308 18392 10310
rect 18416 10308 18472 10310
rect 18496 10308 18552 10310
rect 18256 9274 18312 9276
rect 18336 9274 18392 9276
rect 18416 9274 18472 9276
rect 18496 9274 18552 9276
rect 18256 9222 18282 9274
rect 18282 9222 18312 9274
rect 18336 9222 18346 9274
rect 18346 9222 18392 9274
rect 18416 9222 18462 9274
rect 18462 9222 18472 9274
rect 18496 9222 18526 9274
rect 18526 9222 18552 9274
rect 18256 9220 18312 9222
rect 18336 9220 18392 9222
rect 18416 9220 18472 9222
rect 18496 9220 18552 9222
rect 16756 8730 16812 8732
rect 16836 8730 16892 8732
rect 16916 8730 16972 8732
rect 16996 8730 17052 8732
rect 16756 8678 16782 8730
rect 16782 8678 16812 8730
rect 16836 8678 16846 8730
rect 16846 8678 16892 8730
rect 16916 8678 16962 8730
rect 16962 8678 16972 8730
rect 16996 8678 17026 8730
rect 17026 8678 17052 8730
rect 16756 8676 16812 8678
rect 16836 8676 16892 8678
rect 16916 8676 16972 8678
rect 16996 8676 17052 8678
rect 15256 6010 15312 6012
rect 15336 6010 15392 6012
rect 15416 6010 15472 6012
rect 15496 6010 15552 6012
rect 15256 5958 15282 6010
rect 15282 5958 15312 6010
rect 15336 5958 15346 6010
rect 15346 5958 15392 6010
rect 15416 5958 15462 6010
rect 15462 5958 15472 6010
rect 15496 5958 15526 6010
rect 15526 5958 15552 6010
rect 15256 5956 15312 5958
rect 15336 5956 15392 5958
rect 15416 5956 15472 5958
rect 15496 5956 15552 5958
rect 15256 4922 15312 4924
rect 15336 4922 15392 4924
rect 15416 4922 15472 4924
rect 15496 4922 15552 4924
rect 15256 4870 15282 4922
rect 15282 4870 15312 4922
rect 15336 4870 15346 4922
rect 15346 4870 15392 4922
rect 15416 4870 15462 4922
rect 15462 4870 15472 4922
rect 15496 4870 15526 4922
rect 15526 4870 15552 4922
rect 15256 4868 15312 4870
rect 15336 4868 15392 4870
rect 15416 4868 15472 4870
rect 15496 4868 15552 4870
rect 13756 4378 13812 4380
rect 13836 4378 13892 4380
rect 13916 4378 13972 4380
rect 13996 4378 14052 4380
rect 13756 4326 13782 4378
rect 13782 4326 13812 4378
rect 13836 4326 13846 4378
rect 13846 4326 13892 4378
rect 13916 4326 13962 4378
rect 13962 4326 13972 4378
rect 13996 4326 14026 4378
rect 14026 4326 14052 4378
rect 13756 4324 13812 4326
rect 13836 4324 13892 4326
rect 13916 4324 13972 4326
rect 13996 4324 14052 4326
rect 13756 3290 13812 3292
rect 13836 3290 13892 3292
rect 13916 3290 13972 3292
rect 13996 3290 14052 3292
rect 13756 3238 13782 3290
rect 13782 3238 13812 3290
rect 13836 3238 13846 3290
rect 13846 3238 13892 3290
rect 13916 3238 13962 3290
rect 13962 3238 13972 3290
rect 13996 3238 14026 3290
rect 14026 3238 14052 3290
rect 13756 3236 13812 3238
rect 13836 3236 13892 3238
rect 13916 3236 13972 3238
rect 13996 3236 14052 3238
rect 15256 3834 15312 3836
rect 15336 3834 15392 3836
rect 15416 3834 15472 3836
rect 15496 3834 15552 3836
rect 15256 3782 15282 3834
rect 15282 3782 15312 3834
rect 15336 3782 15346 3834
rect 15346 3782 15392 3834
rect 15416 3782 15462 3834
rect 15462 3782 15472 3834
rect 15496 3782 15526 3834
rect 15526 3782 15552 3834
rect 15256 3780 15312 3782
rect 15336 3780 15392 3782
rect 15416 3780 15472 3782
rect 15496 3780 15552 3782
rect 16756 7642 16812 7644
rect 16836 7642 16892 7644
rect 16916 7642 16972 7644
rect 16996 7642 17052 7644
rect 16756 7590 16782 7642
rect 16782 7590 16812 7642
rect 16836 7590 16846 7642
rect 16846 7590 16892 7642
rect 16916 7590 16962 7642
rect 16962 7590 16972 7642
rect 16996 7590 17026 7642
rect 17026 7590 17052 7642
rect 16756 7588 16812 7590
rect 16836 7588 16892 7590
rect 16916 7588 16972 7590
rect 16996 7588 17052 7590
rect 18256 8186 18312 8188
rect 18336 8186 18392 8188
rect 18416 8186 18472 8188
rect 18496 8186 18552 8188
rect 18256 8134 18282 8186
rect 18282 8134 18312 8186
rect 18336 8134 18346 8186
rect 18346 8134 18392 8186
rect 18416 8134 18462 8186
rect 18462 8134 18472 8186
rect 18496 8134 18526 8186
rect 18526 8134 18552 8186
rect 18256 8132 18312 8134
rect 18336 8132 18392 8134
rect 18416 8132 18472 8134
rect 18496 8132 18552 8134
rect 18256 7098 18312 7100
rect 18336 7098 18392 7100
rect 18416 7098 18472 7100
rect 18496 7098 18552 7100
rect 18256 7046 18282 7098
rect 18282 7046 18312 7098
rect 18336 7046 18346 7098
rect 18346 7046 18392 7098
rect 18416 7046 18462 7098
rect 18462 7046 18472 7098
rect 18496 7046 18526 7098
rect 18526 7046 18552 7098
rect 18256 7044 18312 7046
rect 18336 7044 18392 7046
rect 18416 7044 18472 7046
rect 18496 7044 18552 7046
rect 16756 6554 16812 6556
rect 16836 6554 16892 6556
rect 16916 6554 16972 6556
rect 16996 6554 17052 6556
rect 16756 6502 16782 6554
rect 16782 6502 16812 6554
rect 16836 6502 16846 6554
rect 16846 6502 16892 6554
rect 16916 6502 16962 6554
rect 16962 6502 16972 6554
rect 16996 6502 17026 6554
rect 17026 6502 17052 6554
rect 16756 6500 16812 6502
rect 16836 6500 16892 6502
rect 16916 6500 16972 6502
rect 16996 6500 17052 6502
rect 15256 2746 15312 2748
rect 15336 2746 15392 2748
rect 15416 2746 15472 2748
rect 15496 2746 15552 2748
rect 15256 2694 15282 2746
rect 15282 2694 15312 2746
rect 15336 2694 15346 2746
rect 15346 2694 15392 2746
rect 15416 2694 15462 2746
rect 15462 2694 15472 2746
rect 15496 2694 15526 2746
rect 15526 2694 15552 2746
rect 15256 2692 15312 2694
rect 15336 2692 15392 2694
rect 15416 2692 15472 2694
rect 15496 2692 15552 2694
rect 14370 2488 14426 2544
rect 16756 5466 16812 5468
rect 16836 5466 16892 5468
rect 16916 5466 16972 5468
rect 16996 5466 17052 5468
rect 16756 5414 16782 5466
rect 16782 5414 16812 5466
rect 16836 5414 16846 5466
rect 16846 5414 16892 5466
rect 16916 5414 16962 5466
rect 16962 5414 16972 5466
rect 16996 5414 17026 5466
rect 17026 5414 17052 5466
rect 16756 5412 16812 5414
rect 16836 5412 16892 5414
rect 16916 5412 16972 5414
rect 16996 5412 17052 5414
rect 16756 4378 16812 4380
rect 16836 4378 16892 4380
rect 16916 4378 16972 4380
rect 16996 4378 17052 4380
rect 16756 4326 16782 4378
rect 16782 4326 16812 4378
rect 16836 4326 16846 4378
rect 16846 4326 16892 4378
rect 16916 4326 16962 4378
rect 16962 4326 16972 4378
rect 16996 4326 17026 4378
rect 17026 4326 17052 4378
rect 16756 4324 16812 4326
rect 16836 4324 16892 4326
rect 16916 4324 16972 4326
rect 16996 4324 17052 4326
rect 18256 6010 18312 6012
rect 18336 6010 18392 6012
rect 18416 6010 18472 6012
rect 18496 6010 18552 6012
rect 18256 5958 18282 6010
rect 18282 5958 18312 6010
rect 18336 5958 18346 6010
rect 18346 5958 18392 6010
rect 18416 5958 18462 6010
rect 18462 5958 18472 6010
rect 18496 5958 18526 6010
rect 18526 5958 18552 6010
rect 18256 5956 18312 5958
rect 18336 5956 18392 5958
rect 18416 5956 18472 5958
rect 18496 5956 18552 5958
rect 19756 13082 19812 13084
rect 19836 13082 19892 13084
rect 19916 13082 19972 13084
rect 19996 13082 20052 13084
rect 19756 13030 19782 13082
rect 19782 13030 19812 13082
rect 19836 13030 19846 13082
rect 19846 13030 19892 13082
rect 19916 13030 19962 13082
rect 19962 13030 19972 13082
rect 19996 13030 20026 13082
rect 20026 13030 20052 13082
rect 19756 13028 19812 13030
rect 19836 13028 19892 13030
rect 19916 13028 19972 13030
rect 19996 13028 20052 13030
rect 21256 14714 21312 14716
rect 21336 14714 21392 14716
rect 21416 14714 21472 14716
rect 21496 14714 21552 14716
rect 21256 14662 21282 14714
rect 21282 14662 21312 14714
rect 21336 14662 21346 14714
rect 21346 14662 21392 14714
rect 21416 14662 21462 14714
rect 21462 14662 21472 14714
rect 21496 14662 21526 14714
rect 21526 14662 21552 14714
rect 21256 14660 21312 14662
rect 21336 14660 21392 14662
rect 21416 14660 21472 14662
rect 21496 14660 21552 14662
rect 22756 27226 22812 27228
rect 22836 27226 22892 27228
rect 22916 27226 22972 27228
rect 22996 27226 23052 27228
rect 22756 27174 22782 27226
rect 22782 27174 22812 27226
rect 22836 27174 22846 27226
rect 22846 27174 22892 27226
rect 22916 27174 22962 27226
rect 22962 27174 22972 27226
rect 22996 27174 23026 27226
rect 23026 27174 23052 27226
rect 22756 27172 22812 27174
rect 22836 27172 22892 27174
rect 22916 27172 22972 27174
rect 22996 27172 23052 27174
rect 25756 27226 25812 27228
rect 25836 27226 25892 27228
rect 25916 27226 25972 27228
rect 25996 27226 26052 27228
rect 25756 27174 25782 27226
rect 25782 27174 25812 27226
rect 25836 27174 25846 27226
rect 25846 27174 25892 27226
rect 25916 27174 25962 27226
rect 25962 27174 25972 27226
rect 25996 27174 26026 27226
rect 26026 27174 26052 27226
rect 25756 27172 25812 27174
rect 25836 27172 25892 27174
rect 25916 27172 25972 27174
rect 25996 27172 26052 27174
rect 24256 26682 24312 26684
rect 24336 26682 24392 26684
rect 24416 26682 24472 26684
rect 24496 26682 24552 26684
rect 24256 26630 24282 26682
rect 24282 26630 24312 26682
rect 24336 26630 24346 26682
rect 24346 26630 24392 26682
rect 24416 26630 24462 26682
rect 24462 26630 24472 26682
rect 24496 26630 24526 26682
rect 24526 26630 24552 26682
rect 24256 26628 24312 26630
rect 24336 26628 24392 26630
rect 24416 26628 24472 26630
rect 24496 26628 24552 26630
rect 27256 26682 27312 26684
rect 27336 26682 27392 26684
rect 27416 26682 27472 26684
rect 27496 26682 27552 26684
rect 27256 26630 27282 26682
rect 27282 26630 27312 26682
rect 27336 26630 27346 26682
rect 27346 26630 27392 26682
rect 27416 26630 27462 26682
rect 27462 26630 27472 26682
rect 27496 26630 27526 26682
rect 27526 26630 27552 26682
rect 27256 26628 27312 26630
rect 27336 26628 27392 26630
rect 27416 26628 27472 26630
rect 27496 26628 27552 26630
rect 22756 26138 22812 26140
rect 22836 26138 22892 26140
rect 22916 26138 22972 26140
rect 22996 26138 23052 26140
rect 22756 26086 22782 26138
rect 22782 26086 22812 26138
rect 22836 26086 22846 26138
rect 22846 26086 22892 26138
rect 22916 26086 22962 26138
rect 22962 26086 22972 26138
rect 22996 26086 23026 26138
rect 23026 26086 23052 26138
rect 22756 26084 22812 26086
rect 22836 26084 22892 26086
rect 22916 26084 22972 26086
rect 22996 26084 23052 26086
rect 25756 26138 25812 26140
rect 25836 26138 25892 26140
rect 25916 26138 25972 26140
rect 25996 26138 26052 26140
rect 25756 26086 25782 26138
rect 25782 26086 25812 26138
rect 25836 26086 25846 26138
rect 25846 26086 25892 26138
rect 25916 26086 25962 26138
rect 25962 26086 25972 26138
rect 25996 26086 26026 26138
rect 26026 26086 26052 26138
rect 25756 26084 25812 26086
rect 25836 26084 25892 26086
rect 25916 26084 25972 26086
rect 25996 26084 26052 26086
rect 24256 25594 24312 25596
rect 24336 25594 24392 25596
rect 24416 25594 24472 25596
rect 24496 25594 24552 25596
rect 24256 25542 24282 25594
rect 24282 25542 24312 25594
rect 24336 25542 24346 25594
rect 24346 25542 24392 25594
rect 24416 25542 24462 25594
rect 24462 25542 24472 25594
rect 24496 25542 24526 25594
rect 24526 25542 24552 25594
rect 24256 25540 24312 25542
rect 24336 25540 24392 25542
rect 24416 25540 24472 25542
rect 24496 25540 24552 25542
rect 27256 25594 27312 25596
rect 27336 25594 27392 25596
rect 27416 25594 27472 25596
rect 27496 25594 27552 25596
rect 27256 25542 27282 25594
rect 27282 25542 27312 25594
rect 27336 25542 27346 25594
rect 27346 25542 27392 25594
rect 27416 25542 27462 25594
rect 27462 25542 27472 25594
rect 27496 25542 27526 25594
rect 27526 25542 27552 25594
rect 27256 25540 27312 25542
rect 27336 25540 27392 25542
rect 27416 25540 27472 25542
rect 27496 25540 27552 25542
rect 22756 25050 22812 25052
rect 22836 25050 22892 25052
rect 22916 25050 22972 25052
rect 22996 25050 23052 25052
rect 22756 24998 22782 25050
rect 22782 24998 22812 25050
rect 22836 24998 22846 25050
rect 22846 24998 22892 25050
rect 22916 24998 22962 25050
rect 22962 24998 22972 25050
rect 22996 24998 23026 25050
rect 23026 24998 23052 25050
rect 22756 24996 22812 24998
rect 22836 24996 22892 24998
rect 22916 24996 22972 24998
rect 22996 24996 23052 24998
rect 25756 25050 25812 25052
rect 25836 25050 25892 25052
rect 25916 25050 25972 25052
rect 25996 25050 26052 25052
rect 25756 24998 25782 25050
rect 25782 24998 25812 25050
rect 25836 24998 25846 25050
rect 25846 24998 25892 25050
rect 25916 24998 25962 25050
rect 25962 24998 25972 25050
rect 25996 24998 26026 25050
rect 26026 24998 26052 25050
rect 25756 24996 25812 24998
rect 25836 24996 25892 24998
rect 25916 24996 25972 24998
rect 25996 24996 26052 24998
rect 24256 24506 24312 24508
rect 24336 24506 24392 24508
rect 24416 24506 24472 24508
rect 24496 24506 24552 24508
rect 24256 24454 24282 24506
rect 24282 24454 24312 24506
rect 24336 24454 24346 24506
rect 24346 24454 24392 24506
rect 24416 24454 24462 24506
rect 24462 24454 24472 24506
rect 24496 24454 24526 24506
rect 24526 24454 24552 24506
rect 24256 24452 24312 24454
rect 24336 24452 24392 24454
rect 24416 24452 24472 24454
rect 24496 24452 24552 24454
rect 27256 24506 27312 24508
rect 27336 24506 27392 24508
rect 27416 24506 27472 24508
rect 27496 24506 27552 24508
rect 27256 24454 27282 24506
rect 27282 24454 27312 24506
rect 27336 24454 27346 24506
rect 27346 24454 27392 24506
rect 27416 24454 27462 24506
rect 27462 24454 27472 24506
rect 27496 24454 27526 24506
rect 27526 24454 27552 24506
rect 27256 24452 27312 24454
rect 27336 24452 27392 24454
rect 27416 24452 27472 24454
rect 27496 24452 27552 24454
rect 22756 23962 22812 23964
rect 22836 23962 22892 23964
rect 22916 23962 22972 23964
rect 22996 23962 23052 23964
rect 22756 23910 22782 23962
rect 22782 23910 22812 23962
rect 22836 23910 22846 23962
rect 22846 23910 22892 23962
rect 22916 23910 22962 23962
rect 22962 23910 22972 23962
rect 22996 23910 23026 23962
rect 23026 23910 23052 23962
rect 22756 23908 22812 23910
rect 22836 23908 22892 23910
rect 22916 23908 22972 23910
rect 22996 23908 23052 23910
rect 25756 23962 25812 23964
rect 25836 23962 25892 23964
rect 25916 23962 25972 23964
rect 25996 23962 26052 23964
rect 25756 23910 25782 23962
rect 25782 23910 25812 23962
rect 25836 23910 25846 23962
rect 25846 23910 25892 23962
rect 25916 23910 25962 23962
rect 25962 23910 25972 23962
rect 25996 23910 26026 23962
rect 26026 23910 26052 23962
rect 25756 23908 25812 23910
rect 25836 23908 25892 23910
rect 25916 23908 25972 23910
rect 25996 23908 26052 23910
rect 24256 23418 24312 23420
rect 24336 23418 24392 23420
rect 24416 23418 24472 23420
rect 24496 23418 24552 23420
rect 24256 23366 24282 23418
rect 24282 23366 24312 23418
rect 24336 23366 24346 23418
rect 24346 23366 24392 23418
rect 24416 23366 24462 23418
rect 24462 23366 24472 23418
rect 24496 23366 24526 23418
rect 24526 23366 24552 23418
rect 24256 23364 24312 23366
rect 24336 23364 24392 23366
rect 24416 23364 24472 23366
rect 24496 23364 24552 23366
rect 27256 23418 27312 23420
rect 27336 23418 27392 23420
rect 27416 23418 27472 23420
rect 27496 23418 27552 23420
rect 27256 23366 27282 23418
rect 27282 23366 27312 23418
rect 27336 23366 27346 23418
rect 27346 23366 27392 23418
rect 27416 23366 27462 23418
rect 27462 23366 27472 23418
rect 27496 23366 27526 23418
rect 27526 23366 27552 23418
rect 27256 23364 27312 23366
rect 27336 23364 27392 23366
rect 27416 23364 27472 23366
rect 27496 23364 27552 23366
rect 22756 22874 22812 22876
rect 22836 22874 22892 22876
rect 22916 22874 22972 22876
rect 22996 22874 23052 22876
rect 22756 22822 22782 22874
rect 22782 22822 22812 22874
rect 22836 22822 22846 22874
rect 22846 22822 22892 22874
rect 22916 22822 22962 22874
rect 22962 22822 22972 22874
rect 22996 22822 23026 22874
rect 23026 22822 23052 22874
rect 22756 22820 22812 22822
rect 22836 22820 22892 22822
rect 22916 22820 22972 22822
rect 22996 22820 23052 22822
rect 25756 22874 25812 22876
rect 25836 22874 25892 22876
rect 25916 22874 25972 22876
rect 25996 22874 26052 22876
rect 25756 22822 25782 22874
rect 25782 22822 25812 22874
rect 25836 22822 25846 22874
rect 25846 22822 25892 22874
rect 25916 22822 25962 22874
rect 25962 22822 25972 22874
rect 25996 22822 26026 22874
rect 26026 22822 26052 22874
rect 25756 22820 25812 22822
rect 25836 22820 25892 22822
rect 25916 22820 25972 22822
rect 25996 22820 26052 22822
rect 24256 22330 24312 22332
rect 24336 22330 24392 22332
rect 24416 22330 24472 22332
rect 24496 22330 24552 22332
rect 24256 22278 24282 22330
rect 24282 22278 24312 22330
rect 24336 22278 24346 22330
rect 24346 22278 24392 22330
rect 24416 22278 24462 22330
rect 24462 22278 24472 22330
rect 24496 22278 24526 22330
rect 24526 22278 24552 22330
rect 24256 22276 24312 22278
rect 24336 22276 24392 22278
rect 24416 22276 24472 22278
rect 24496 22276 24552 22278
rect 27256 22330 27312 22332
rect 27336 22330 27392 22332
rect 27416 22330 27472 22332
rect 27496 22330 27552 22332
rect 27256 22278 27282 22330
rect 27282 22278 27312 22330
rect 27336 22278 27346 22330
rect 27346 22278 27392 22330
rect 27416 22278 27462 22330
rect 27462 22278 27472 22330
rect 27496 22278 27526 22330
rect 27526 22278 27552 22330
rect 27256 22276 27312 22278
rect 27336 22276 27392 22278
rect 27416 22276 27472 22278
rect 27496 22276 27552 22278
rect 22756 21786 22812 21788
rect 22836 21786 22892 21788
rect 22916 21786 22972 21788
rect 22996 21786 23052 21788
rect 22756 21734 22782 21786
rect 22782 21734 22812 21786
rect 22836 21734 22846 21786
rect 22846 21734 22892 21786
rect 22916 21734 22962 21786
rect 22962 21734 22972 21786
rect 22996 21734 23026 21786
rect 23026 21734 23052 21786
rect 22756 21732 22812 21734
rect 22836 21732 22892 21734
rect 22916 21732 22972 21734
rect 22996 21732 23052 21734
rect 25756 21786 25812 21788
rect 25836 21786 25892 21788
rect 25916 21786 25972 21788
rect 25996 21786 26052 21788
rect 25756 21734 25782 21786
rect 25782 21734 25812 21786
rect 25836 21734 25846 21786
rect 25846 21734 25892 21786
rect 25916 21734 25962 21786
rect 25962 21734 25972 21786
rect 25996 21734 26026 21786
rect 26026 21734 26052 21786
rect 25756 21732 25812 21734
rect 25836 21732 25892 21734
rect 25916 21732 25972 21734
rect 25996 21732 26052 21734
rect 24256 21242 24312 21244
rect 24336 21242 24392 21244
rect 24416 21242 24472 21244
rect 24496 21242 24552 21244
rect 24256 21190 24282 21242
rect 24282 21190 24312 21242
rect 24336 21190 24346 21242
rect 24346 21190 24392 21242
rect 24416 21190 24462 21242
rect 24462 21190 24472 21242
rect 24496 21190 24526 21242
rect 24526 21190 24552 21242
rect 24256 21188 24312 21190
rect 24336 21188 24392 21190
rect 24416 21188 24472 21190
rect 24496 21188 24552 21190
rect 27256 21242 27312 21244
rect 27336 21242 27392 21244
rect 27416 21242 27472 21244
rect 27496 21242 27552 21244
rect 27256 21190 27282 21242
rect 27282 21190 27312 21242
rect 27336 21190 27346 21242
rect 27346 21190 27392 21242
rect 27416 21190 27462 21242
rect 27462 21190 27472 21242
rect 27496 21190 27526 21242
rect 27526 21190 27552 21242
rect 27256 21188 27312 21190
rect 27336 21188 27392 21190
rect 27416 21188 27472 21190
rect 27496 21188 27552 21190
rect 22756 20698 22812 20700
rect 22836 20698 22892 20700
rect 22916 20698 22972 20700
rect 22996 20698 23052 20700
rect 22756 20646 22782 20698
rect 22782 20646 22812 20698
rect 22836 20646 22846 20698
rect 22846 20646 22892 20698
rect 22916 20646 22962 20698
rect 22962 20646 22972 20698
rect 22996 20646 23026 20698
rect 23026 20646 23052 20698
rect 22756 20644 22812 20646
rect 22836 20644 22892 20646
rect 22916 20644 22972 20646
rect 22996 20644 23052 20646
rect 25756 20698 25812 20700
rect 25836 20698 25892 20700
rect 25916 20698 25972 20700
rect 25996 20698 26052 20700
rect 25756 20646 25782 20698
rect 25782 20646 25812 20698
rect 25836 20646 25846 20698
rect 25846 20646 25892 20698
rect 25916 20646 25962 20698
rect 25962 20646 25972 20698
rect 25996 20646 26026 20698
rect 26026 20646 26052 20698
rect 25756 20644 25812 20646
rect 25836 20644 25892 20646
rect 25916 20644 25972 20646
rect 25996 20644 26052 20646
rect 24256 20154 24312 20156
rect 24336 20154 24392 20156
rect 24416 20154 24472 20156
rect 24496 20154 24552 20156
rect 24256 20102 24282 20154
rect 24282 20102 24312 20154
rect 24336 20102 24346 20154
rect 24346 20102 24392 20154
rect 24416 20102 24462 20154
rect 24462 20102 24472 20154
rect 24496 20102 24526 20154
rect 24526 20102 24552 20154
rect 24256 20100 24312 20102
rect 24336 20100 24392 20102
rect 24416 20100 24472 20102
rect 24496 20100 24552 20102
rect 27256 20154 27312 20156
rect 27336 20154 27392 20156
rect 27416 20154 27472 20156
rect 27496 20154 27552 20156
rect 27256 20102 27282 20154
rect 27282 20102 27312 20154
rect 27336 20102 27346 20154
rect 27346 20102 27392 20154
rect 27416 20102 27462 20154
rect 27462 20102 27472 20154
rect 27496 20102 27526 20154
rect 27526 20102 27552 20154
rect 27256 20100 27312 20102
rect 27336 20100 27392 20102
rect 27416 20100 27472 20102
rect 27496 20100 27552 20102
rect 22756 19610 22812 19612
rect 22836 19610 22892 19612
rect 22916 19610 22972 19612
rect 22996 19610 23052 19612
rect 22756 19558 22782 19610
rect 22782 19558 22812 19610
rect 22836 19558 22846 19610
rect 22846 19558 22892 19610
rect 22916 19558 22962 19610
rect 22962 19558 22972 19610
rect 22996 19558 23026 19610
rect 23026 19558 23052 19610
rect 22756 19556 22812 19558
rect 22836 19556 22892 19558
rect 22916 19556 22972 19558
rect 22996 19556 23052 19558
rect 25756 19610 25812 19612
rect 25836 19610 25892 19612
rect 25916 19610 25972 19612
rect 25996 19610 26052 19612
rect 25756 19558 25782 19610
rect 25782 19558 25812 19610
rect 25836 19558 25846 19610
rect 25846 19558 25892 19610
rect 25916 19558 25962 19610
rect 25962 19558 25972 19610
rect 25996 19558 26026 19610
rect 26026 19558 26052 19610
rect 25756 19556 25812 19558
rect 25836 19556 25892 19558
rect 25916 19556 25972 19558
rect 25996 19556 26052 19558
rect 24256 19066 24312 19068
rect 24336 19066 24392 19068
rect 24416 19066 24472 19068
rect 24496 19066 24552 19068
rect 24256 19014 24282 19066
rect 24282 19014 24312 19066
rect 24336 19014 24346 19066
rect 24346 19014 24392 19066
rect 24416 19014 24462 19066
rect 24462 19014 24472 19066
rect 24496 19014 24526 19066
rect 24526 19014 24552 19066
rect 24256 19012 24312 19014
rect 24336 19012 24392 19014
rect 24416 19012 24472 19014
rect 24496 19012 24552 19014
rect 27256 19066 27312 19068
rect 27336 19066 27392 19068
rect 27416 19066 27472 19068
rect 27496 19066 27552 19068
rect 27256 19014 27282 19066
rect 27282 19014 27312 19066
rect 27336 19014 27346 19066
rect 27346 19014 27392 19066
rect 27416 19014 27462 19066
rect 27462 19014 27472 19066
rect 27496 19014 27526 19066
rect 27526 19014 27552 19066
rect 27256 19012 27312 19014
rect 27336 19012 27392 19014
rect 27416 19012 27472 19014
rect 27496 19012 27552 19014
rect 22756 18522 22812 18524
rect 22836 18522 22892 18524
rect 22916 18522 22972 18524
rect 22996 18522 23052 18524
rect 22756 18470 22782 18522
rect 22782 18470 22812 18522
rect 22836 18470 22846 18522
rect 22846 18470 22892 18522
rect 22916 18470 22962 18522
rect 22962 18470 22972 18522
rect 22996 18470 23026 18522
rect 23026 18470 23052 18522
rect 22756 18468 22812 18470
rect 22836 18468 22892 18470
rect 22916 18468 22972 18470
rect 22996 18468 23052 18470
rect 25756 18522 25812 18524
rect 25836 18522 25892 18524
rect 25916 18522 25972 18524
rect 25996 18522 26052 18524
rect 25756 18470 25782 18522
rect 25782 18470 25812 18522
rect 25836 18470 25846 18522
rect 25846 18470 25892 18522
rect 25916 18470 25962 18522
rect 25962 18470 25972 18522
rect 25996 18470 26026 18522
rect 26026 18470 26052 18522
rect 25756 18468 25812 18470
rect 25836 18468 25892 18470
rect 25916 18468 25972 18470
rect 25996 18468 26052 18470
rect 24256 17978 24312 17980
rect 24336 17978 24392 17980
rect 24416 17978 24472 17980
rect 24496 17978 24552 17980
rect 24256 17926 24282 17978
rect 24282 17926 24312 17978
rect 24336 17926 24346 17978
rect 24346 17926 24392 17978
rect 24416 17926 24462 17978
rect 24462 17926 24472 17978
rect 24496 17926 24526 17978
rect 24526 17926 24552 17978
rect 24256 17924 24312 17926
rect 24336 17924 24392 17926
rect 24416 17924 24472 17926
rect 24496 17924 24552 17926
rect 27256 17978 27312 17980
rect 27336 17978 27392 17980
rect 27416 17978 27472 17980
rect 27496 17978 27552 17980
rect 27256 17926 27282 17978
rect 27282 17926 27312 17978
rect 27336 17926 27346 17978
rect 27346 17926 27392 17978
rect 27416 17926 27462 17978
rect 27462 17926 27472 17978
rect 27496 17926 27526 17978
rect 27526 17926 27552 17978
rect 27256 17924 27312 17926
rect 27336 17924 27392 17926
rect 27416 17924 27472 17926
rect 27496 17924 27552 17926
rect 22756 17434 22812 17436
rect 22836 17434 22892 17436
rect 22916 17434 22972 17436
rect 22996 17434 23052 17436
rect 22756 17382 22782 17434
rect 22782 17382 22812 17434
rect 22836 17382 22846 17434
rect 22846 17382 22892 17434
rect 22916 17382 22962 17434
rect 22962 17382 22972 17434
rect 22996 17382 23026 17434
rect 23026 17382 23052 17434
rect 22756 17380 22812 17382
rect 22836 17380 22892 17382
rect 22916 17380 22972 17382
rect 22996 17380 23052 17382
rect 25756 17434 25812 17436
rect 25836 17434 25892 17436
rect 25916 17434 25972 17436
rect 25996 17434 26052 17436
rect 25756 17382 25782 17434
rect 25782 17382 25812 17434
rect 25836 17382 25846 17434
rect 25846 17382 25892 17434
rect 25916 17382 25962 17434
rect 25962 17382 25972 17434
rect 25996 17382 26026 17434
rect 26026 17382 26052 17434
rect 25756 17380 25812 17382
rect 25836 17380 25892 17382
rect 25916 17380 25972 17382
rect 25996 17380 26052 17382
rect 24256 16890 24312 16892
rect 24336 16890 24392 16892
rect 24416 16890 24472 16892
rect 24496 16890 24552 16892
rect 24256 16838 24282 16890
rect 24282 16838 24312 16890
rect 24336 16838 24346 16890
rect 24346 16838 24392 16890
rect 24416 16838 24462 16890
rect 24462 16838 24472 16890
rect 24496 16838 24526 16890
rect 24526 16838 24552 16890
rect 24256 16836 24312 16838
rect 24336 16836 24392 16838
rect 24416 16836 24472 16838
rect 24496 16836 24552 16838
rect 27256 16890 27312 16892
rect 27336 16890 27392 16892
rect 27416 16890 27472 16892
rect 27496 16890 27552 16892
rect 27256 16838 27282 16890
rect 27282 16838 27312 16890
rect 27336 16838 27346 16890
rect 27346 16838 27392 16890
rect 27416 16838 27462 16890
rect 27462 16838 27472 16890
rect 27496 16838 27526 16890
rect 27526 16838 27552 16890
rect 27256 16836 27312 16838
rect 27336 16836 27392 16838
rect 27416 16836 27472 16838
rect 27496 16836 27552 16838
rect 22756 16346 22812 16348
rect 22836 16346 22892 16348
rect 22916 16346 22972 16348
rect 22996 16346 23052 16348
rect 22756 16294 22782 16346
rect 22782 16294 22812 16346
rect 22836 16294 22846 16346
rect 22846 16294 22892 16346
rect 22916 16294 22962 16346
rect 22962 16294 22972 16346
rect 22996 16294 23026 16346
rect 23026 16294 23052 16346
rect 22756 16292 22812 16294
rect 22836 16292 22892 16294
rect 22916 16292 22972 16294
rect 22996 16292 23052 16294
rect 25756 16346 25812 16348
rect 25836 16346 25892 16348
rect 25916 16346 25972 16348
rect 25996 16346 26052 16348
rect 25756 16294 25782 16346
rect 25782 16294 25812 16346
rect 25836 16294 25846 16346
rect 25846 16294 25892 16346
rect 25916 16294 25962 16346
rect 25962 16294 25972 16346
rect 25996 16294 26026 16346
rect 26026 16294 26052 16346
rect 25756 16292 25812 16294
rect 25836 16292 25892 16294
rect 25916 16292 25972 16294
rect 25996 16292 26052 16294
rect 24256 15802 24312 15804
rect 24336 15802 24392 15804
rect 24416 15802 24472 15804
rect 24496 15802 24552 15804
rect 24256 15750 24282 15802
rect 24282 15750 24312 15802
rect 24336 15750 24346 15802
rect 24346 15750 24392 15802
rect 24416 15750 24462 15802
rect 24462 15750 24472 15802
rect 24496 15750 24526 15802
rect 24526 15750 24552 15802
rect 24256 15748 24312 15750
rect 24336 15748 24392 15750
rect 24416 15748 24472 15750
rect 24496 15748 24552 15750
rect 27256 15802 27312 15804
rect 27336 15802 27392 15804
rect 27416 15802 27472 15804
rect 27496 15802 27552 15804
rect 27256 15750 27282 15802
rect 27282 15750 27312 15802
rect 27336 15750 27346 15802
rect 27346 15750 27392 15802
rect 27416 15750 27462 15802
rect 27462 15750 27472 15802
rect 27496 15750 27526 15802
rect 27526 15750 27552 15802
rect 27256 15748 27312 15750
rect 27336 15748 27392 15750
rect 27416 15748 27472 15750
rect 27496 15748 27552 15750
rect 22756 15258 22812 15260
rect 22836 15258 22892 15260
rect 22916 15258 22972 15260
rect 22996 15258 23052 15260
rect 22756 15206 22782 15258
rect 22782 15206 22812 15258
rect 22836 15206 22846 15258
rect 22846 15206 22892 15258
rect 22916 15206 22962 15258
rect 22962 15206 22972 15258
rect 22996 15206 23026 15258
rect 23026 15206 23052 15258
rect 22756 15204 22812 15206
rect 22836 15204 22892 15206
rect 22916 15204 22972 15206
rect 22996 15204 23052 15206
rect 25756 15258 25812 15260
rect 25836 15258 25892 15260
rect 25916 15258 25972 15260
rect 25996 15258 26052 15260
rect 25756 15206 25782 15258
rect 25782 15206 25812 15258
rect 25836 15206 25846 15258
rect 25846 15206 25892 15258
rect 25916 15206 25962 15258
rect 25962 15206 25972 15258
rect 25996 15206 26026 15258
rect 26026 15206 26052 15258
rect 25756 15204 25812 15206
rect 25836 15204 25892 15206
rect 25916 15204 25972 15206
rect 25996 15204 26052 15206
rect 24256 14714 24312 14716
rect 24336 14714 24392 14716
rect 24416 14714 24472 14716
rect 24496 14714 24552 14716
rect 24256 14662 24282 14714
rect 24282 14662 24312 14714
rect 24336 14662 24346 14714
rect 24346 14662 24392 14714
rect 24416 14662 24462 14714
rect 24462 14662 24472 14714
rect 24496 14662 24526 14714
rect 24526 14662 24552 14714
rect 24256 14660 24312 14662
rect 24336 14660 24392 14662
rect 24416 14660 24472 14662
rect 24496 14660 24552 14662
rect 27256 14714 27312 14716
rect 27336 14714 27392 14716
rect 27416 14714 27472 14716
rect 27496 14714 27552 14716
rect 27256 14662 27282 14714
rect 27282 14662 27312 14714
rect 27336 14662 27346 14714
rect 27346 14662 27392 14714
rect 27416 14662 27462 14714
rect 27462 14662 27472 14714
rect 27496 14662 27526 14714
rect 27526 14662 27552 14714
rect 27256 14660 27312 14662
rect 27336 14660 27392 14662
rect 27416 14660 27472 14662
rect 27496 14660 27552 14662
rect 22756 14170 22812 14172
rect 22836 14170 22892 14172
rect 22916 14170 22972 14172
rect 22996 14170 23052 14172
rect 22756 14118 22782 14170
rect 22782 14118 22812 14170
rect 22836 14118 22846 14170
rect 22846 14118 22892 14170
rect 22916 14118 22962 14170
rect 22962 14118 22972 14170
rect 22996 14118 23026 14170
rect 23026 14118 23052 14170
rect 22756 14116 22812 14118
rect 22836 14116 22892 14118
rect 22916 14116 22972 14118
rect 22996 14116 23052 14118
rect 25756 14170 25812 14172
rect 25836 14170 25892 14172
rect 25916 14170 25972 14172
rect 25996 14170 26052 14172
rect 25756 14118 25782 14170
rect 25782 14118 25812 14170
rect 25836 14118 25846 14170
rect 25846 14118 25892 14170
rect 25916 14118 25962 14170
rect 25962 14118 25972 14170
rect 25996 14118 26026 14170
rect 26026 14118 26052 14170
rect 25756 14116 25812 14118
rect 25836 14116 25892 14118
rect 25916 14116 25972 14118
rect 25996 14116 26052 14118
rect 21256 13626 21312 13628
rect 21336 13626 21392 13628
rect 21416 13626 21472 13628
rect 21496 13626 21552 13628
rect 21256 13574 21282 13626
rect 21282 13574 21312 13626
rect 21336 13574 21346 13626
rect 21346 13574 21392 13626
rect 21416 13574 21462 13626
rect 21462 13574 21472 13626
rect 21496 13574 21526 13626
rect 21526 13574 21552 13626
rect 21256 13572 21312 13574
rect 21336 13572 21392 13574
rect 21416 13572 21472 13574
rect 21496 13572 21552 13574
rect 19338 11736 19394 11792
rect 19756 11994 19812 11996
rect 19836 11994 19892 11996
rect 19916 11994 19972 11996
rect 19996 11994 20052 11996
rect 19756 11942 19782 11994
rect 19782 11942 19812 11994
rect 19836 11942 19846 11994
rect 19846 11942 19892 11994
rect 19916 11942 19962 11994
rect 19962 11942 19972 11994
rect 19996 11942 20026 11994
rect 20026 11942 20052 11994
rect 19756 11940 19812 11942
rect 19836 11940 19892 11942
rect 19916 11940 19972 11942
rect 19996 11940 20052 11942
rect 21256 12538 21312 12540
rect 21336 12538 21392 12540
rect 21416 12538 21472 12540
rect 21496 12538 21552 12540
rect 21256 12486 21282 12538
rect 21282 12486 21312 12538
rect 21336 12486 21346 12538
rect 21346 12486 21392 12538
rect 21416 12486 21462 12538
rect 21462 12486 21472 12538
rect 21496 12486 21526 12538
rect 21526 12486 21552 12538
rect 21256 12484 21312 12486
rect 21336 12484 21392 12486
rect 21416 12484 21472 12486
rect 21496 12484 21552 12486
rect 19756 10906 19812 10908
rect 19836 10906 19892 10908
rect 19916 10906 19972 10908
rect 19996 10906 20052 10908
rect 19756 10854 19782 10906
rect 19782 10854 19812 10906
rect 19836 10854 19846 10906
rect 19846 10854 19892 10906
rect 19916 10854 19962 10906
rect 19962 10854 19972 10906
rect 19996 10854 20026 10906
rect 20026 10854 20052 10906
rect 19756 10852 19812 10854
rect 19836 10852 19892 10854
rect 19916 10852 19972 10854
rect 19996 10852 20052 10854
rect 21256 11450 21312 11452
rect 21336 11450 21392 11452
rect 21416 11450 21472 11452
rect 21496 11450 21552 11452
rect 21256 11398 21282 11450
rect 21282 11398 21312 11450
rect 21336 11398 21346 11450
rect 21346 11398 21392 11450
rect 21416 11398 21462 11450
rect 21462 11398 21472 11450
rect 21496 11398 21526 11450
rect 21526 11398 21552 11450
rect 21256 11396 21312 11398
rect 21336 11396 21392 11398
rect 21416 11396 21472 11398
rect 21496 11396 21552 11398
rect 24256 13626 24312 13628
rect 24336 13626 24392 13628
rect 24416 13626 24472 13628
rect 24496 13626 24552 13628
rect 24256 13574 24282 13626
rect 24282 13574 24312 13626
rect 24336 13574 24346 13626
rect 24346 13574 24392 13626
rect 24416 13574 24462 13626
rect 24462 13574 24472 13626
rect 24496 13574 24526 13626
rect 24526 13574 24552 13626
rect 24256 13572 24312 13574
rect 24336 13572 24392 13574
rect 24416 13572 24472 13574
rect 24496 13572 24552 13574
rect 27256 13626 27312 13628
rect 27336 13626 27392 13628
rect 27416 13626 27472 13628
rect 27496 13626 27552 13628
rect 27256 13574 27282 13626
rect 27282 13574 27312 13626
rect 27336 13574 27346 13626
rect 27346 13574 27392 13626
rect 27416 13574 27462 13626
rect 27462 13574 27472 13626
rect 27496 13574 27526 13626
rect 27526 13574 27552 13626
rect 27256 13572 27312 13574
rect 27336 13572 27392 13574
rect 27416 13572 27472 13574
rect 27496 13572 27552 13574
rect 22756 13082 22812 13084
rect 22836 13082 22892 13084
rect 22916 13082 22972 13084
rect 22996 13082 23052 13084
rect 22756 13030 22782 13082
rect 22782 13030 22812 13082
rect 22836 13030 22846 13082
rect 22846 13030 22892 13082
rect 22916 13030 22962 13082
rect 22962 13030 22972 13082
rect 22996 13030 23026 13082
rect 23026 13030 23052 13082
rect 22756 13028 22812 13030
rect 22836 13028 22892 13030
rect 22916 13028 22972 13030
rect 22996 13028 23052 13030
rect 25756 13082 25812 13084
rect 25836 13082 25892 13084
rect 25916 13082 25972 13084
rect 25996 13082 26052 13084
rect 25756 13030 25782 13082
rect 25782 13030 25812 13082
rect 25836 13030 25846 13082
rect 25846 13030 25892 13082
rect 25916 13030 25962 13082
rect 25962 13030 25972 13082
rect 25996 13030 26026 13082
rect 26026 13030 26052 13082
rect 25756 13028 25812 13030
rect 25836 13028 25892 13030
rect 25916 13028 25972 13030
rect 25996 13028 26052 13030
rect 24256 12538 24312 12540
rect 24336 12538 24392 12540
rect 24416 12538 24472 12540
rect 24496 12538 24552 12540
rect 24256 12486 24282 12538
rect 24282 12486 24312 12538
rect 24336 12486 24346 12538
rect 24346 12486 24392 12538
rect 24416 12486 24462 12538
rect 24462 12486 24472 12538
rect 24496 12486 24526 12538
rect 24526 12486 24552 12538
rect 24256 12484 24312 12486
rect 24336 12484 24392 12486
rect 24416 12484 24472 12486
rect 24496 12484 24552 12486
rect 27256 12538 27312 12540
rect 27336 12538 27392 12540
rect 27416 12538 27472 12540
rect 27496 12538 27552 12540
rect 27256 12486 27282 12538
rect 27282 12486 27312 12538
rect 27336 12486 27346 12538
rect 27346 12486 27392 12538
rect 27416 12486 27462 12538
rect 27462 12486 27472 12538
rect 27496 12486 27526 12538
rect 27526 12486 27552 12538
rect 27256 12484 27312 12486
rect 27336 12484 27392 12486
rect 27416 12484 27472 12486
rect 27496 12484 27552 12486
rect 23478 12144 23534 12200
rect 22756 11994 22812 11996
rect 22836 11994 22892 11996
rect 22916 11994 22972 11996
rect 22996 11994 23052 11996
rect 22756 11942 22782 11994
rect 22782 11942 22812 11994
rect 22836 11942 22846 11994
rect 22846 11942 22892 11994
rect 22916 11942 22962 11994
rect 22962 11942 22972 11994
rect 22996 11942 23026 11994
rect 23026 11942 23052 11994
rect 25756 11994 25812 11996
rect 25836 11994 25892 11996
rect 25916 11994 25972 11996
rect 25996 11994 26052 11996
rect 22756 11940 22812 11942
rect 22836 11940 22892 11942
rect 22916 11940 22972 11942
rect 22996 11940 23052 11942
rect 25756 11942 25782 11994
rect 25782 11942 25812 11994
rect 25836 11942 25846 11994
rect 25846 11942 25892 11994
rect 25916 11942 25962 11994
rect 25962 11942 25972 11994
rect 25996 11942 26026 11994
rect 26026 11942 26052 11994
rect 25756 11940 25812 11942
rect 25836 11940 25892 11942
rect 25916 11940 25972 11942
rect 25996 11940 26052 11942
rect 24256 11450 24312 11452
rect 24336 11450 24392 11452
rect 24416 11450 24472 11452
rect 24496 11450 24552 11452
rect 24256 11398 24282 11450
rect 24282 11398 24312 11450
rect 24336 11398 24346 11450
rect 24346 11398 24392 11450
rect 24416 11398 24462 11450
rect 24462 11398 24472 11450
rect 24496 11398 24526 11450
rect 24526 11398 24552 11450
rect 24256 11396 24312 11398
rect 24336 11396 24392 11398
rect 24416 11396 24472 11398
rect 24496 11396 24552 11398
rect 27256 11450 27312 11452
rect 27336 11450 27392 11452
rect 27416 11450 27472 11452
rect 27496 11450 27552 11452
rect 27256 11398 27282 11450
rect 27282 11398 27312 11450
rect 27336 11398 27346 11450
rect 27346 11398 27392 11450
rect 27416 11398 27462 11450
rect 27462 11398 27472 11450
rect 27496 11398 27526 11450
rect 27526 11398 27552 11450
rect 27256 11396 27312 11398
rect 27336 11396 27392 11398
rect 27416 11396 27472 11398
rect 27496 11396 27552 11398
rect 28722 11056 28778 11112
rect 21256 10362 21312 10364
rect 21336 10362 21392 10364
rect 21416 10362 21472 10364
rect 21496 10362 21552 10364
rect 21256 10310 21282 10362
rect 21282 10310 21312 10362
rect 21336 10310 21346 10362
rect 21346 10310 21392 10362
rect 21416 10310 21462 10362
rect 21462 10310 21472 10362
rect 21496 10310 21526 10362
rect 21526 10310 21552 10362
rect 21256 10308 21312 10310
rect 21336 10308 21392 10310
rect 21416 10308 21472 10310
rect 21496 10308 21552 10310
rect 19756 9818 19812 9820
rect 19836 9818 19892 9820
rect 19916 9818 19972 9820
rect 19996 9818 20052 9820
rect 19756 9766 19782 9818
rect 19782 9766 19812 9818
rect 19836 9766 19846 9818
rect 19846 9766 19892 9818
rect 19916 9766 19962 9818
rect 19962 9766 19972 9818
rect 19996 9766 20026 9818
rect 20026 9766 20052 9818
rect 19756 9764 19812 9766
rect 19836 9764 19892 9766
rect 19916 9764 19972 9766
rect 19996 9764 20052 9766
rect 19756 8730 19812 8732
rect 19836 8730 19892 8732
rect 19916 8730 19972 8732
rect 19996 8730 20052 8732
rect 19756 8678 19782 8730
rect 19782 8678 19812 8730
rect 19836 8678 19846 8730
rect 19846 8678 19892 8730
rect 19916 8678 19962 8730
rect 19962 8678 19972 8730
rect 19996 8678 20026 8730
rect 20026 8678 20052 8730
rect 19756 8676 19812 8678
rect 19836 8676 19892 8678
rect 19916 8676 19972 8678
rect 19996 8676 20052 8678
rect 21256 9274 21312 9276
rect 21336 9274 21392 9276
rect 21416 9274 21472 9276
rect 21496 9274 21552 9276
rect 21256 9222 21282 9274
rect 21282 9222 21312 9274
rect 21336 9222 21346 9274
rect 21346 9222 21392 9274
rect 21416 9222 21462 9274
rect 21462 9222 21472 9274
rect 21496 9222 21526 9274
rect 21526 9222 21552 9274
rect 21256 9220 21312 9222
rect 21336 9220 21392 9222
rect 21416 9220 21472 9222
rect 21496 9220 21552 9222
rect 19756 7642 19812 7644
rect 19836 7642 19892 7644
rect 19916 7642 19972 7644
rect 19996 7642 20052 7644
rect 19756 7590 19782 7642
rect 19782 7590 19812 7642
rect 19836 7590 19846 7642
rect 19846 7590 19892 7642
rect 19916 7590 19962 7642
rect 19962 7590 19972 7642
rect 19996 7590 20026 7642
rect 20026 7590 20052 7642
rect 19756 7588 19812 7590
rect 19836 7588 19892 7590
rect 19916 7588 19972 7590
rect 19996 7588 20052 7590
rect 19756 6554 19812 6556
rect 19836 6554 19892 6556
rect 19916 6554 19972 6556
rect 19996 6554 20052 6556
rect 19756 6502 19782 6554
rect 19782 6502 19812 6554
rect 19836 6502 19846 6554
rect 19846 6502 19892 6554
rect 19916 6502 19962 6554
rect 19962 6502 19972 6554
rect 19996 6502 20026 6554
rect 20026 6502 20052 6554
rect 19756 6500 19812 6502
rect 19836 6500 19892 6502
rect 19916 6500 19972 6502
rect 19996 6500 20052 6502
rect 21256 8186 21312 8188
rect 21336 8186 21392 8188
rect 21416 8186 21472 8188
rect 21496 8186 21552 8188
rect 21256 8134 21282 8186
rect 21282 8134 21312 8186
rect 21336 8134 21346 8186
rect 21346 8134 21392 8186
rect 21416 8134 21462 8186
rect 21462 8134 21472 8186
rect 21496 8134 21526 8186
rect 21526 8134 21552 8186
rect 21256 8132 21312 8134
rect 21336 8132 21392 8134
rect 21416 8132 21472 8134
rect 21496 8132 21552 8134
rect 22756 10906 22812 10908
rect 22836 10906 22892 10908
rect 22916 10906 22972 10908
rect 22996 10906 23052 10908
rect 22756 10854 22782 10906
rect 22782 10854 22812 10906
rect 22836 10854 22846 10906
rect 22846 10854 22892 10906
rect 22916 10854 22962 10906
rect 22962 10854 22972 10906
rect 22996 10854 23026 10906
rect 23026 10854 23052 10906
rect 22756 10852 22812 10854
rect 22836 10852 22892 10854
rect 22916 10852 22972 10854
rect 22996 10852 23052 10854
rect 25756 10906 25812 10908
rect 25836 10906 25892 10908
rect 25916 10906 25972 10908
rect 25996 10906 26052 10908
rect 25756 10854 25782 10906
rect 25782 10854 25812 10906
rect 25836 10854 25846 10906
rect 25846 10854 25892 10906
rect 25916 10854 25962 10906
rect 25962 10854 25972 10906
rect 25996 10854 26026 10906
rect 26026 10854 26052 10906
rect 25756 10852 25812 10854
rect 25836 10852 25892 10854
rect 25916 10852 25972 10854
rect 25996 10852 26052 10854
rect 21256 7098 21312 7100
rect 21336 7098 21392 7100
rect 21416 7098 21472 7100
rect 21496 7098 21552 7100
rect 21256 7046 21282 7098
rect 21282 7046 21312 7098
rect 21336 7046 21346 7098
rect 21346 7046 21392 7098
rect 21416 7046 21462 7098
rect 21462 7046 21472 7098
rect 21496 7046 21526 7098
rect 21526 7046 21552 7098
rect 21256 7044 21312 7046
rect 21336 7044 21392 7046
rect 21416 7044 21472 7046
rect 21496 7044 21552 7046
rect 19756 5466 19812 5468
rect 19836 5466 19892 5468
rect 19916 5466 19972 5468
rect 19996 5466 20052 5468
rect 19756 5414 19782 5466
rect 19782 5414 19812 5466
rect 19836 5414 19846 5466
rect 19846 5414 19892 5466
rect 19916 5414 19962 5466
rect 19962 5414 19972 5466
rect 19996 5414 20026 5466
rect 20026 5414 20052 5466
rect 19756 5412 19812 5414
rect 19836 5412 19892 5414
rect 19916 5412 19972 5414
rect 19996 5412 20052 5414
rect 18256 4922 18312 4924
rect 18336 4922 18392 4924
rect 18416 4922 18472 4924
rect 18496 4922 18552 4924
rect 18256 4870 18282 4922
rect 18282 4870 18312 4922
rect 18336 4870 18346 4922
rect 18346 4870 18392 4922
rect 18416 4870 18462 4922
rect 18462 4870 18472 4922
rect 18496 4870 18526 4922
rect 18526 4870 18552 4922
rect 18256 4868 18312 4870
rect 18336 4868 18392 4870
rect 18416 4868 18472 4870
rect 18496 4868 18552 4870
rect 18256 3834 18312 3836
rect 18336 3834 18392 3836
rect 18416 3834 18472 3836
rect 18496 3834 18552 3836
rect 18256 3782 18282 3834
rect 18282 3782 18312 3834
rect 18336 3782 18346 3834
rect 18346 3782 18392 3834
rect 18416 3782 18462 3834
rect 18462 3782 18472 3834
rect 18496 3782 18526 3834
rect 18526 3782 18552 3834
rect 18256 3780 18312 3782
rect 18336 3780 18392 3782
rect 18416 3780 18472 3782
rect 18496 3780 18552 3782
rect 16756 3290 16812 3292
rect 16836 3290 16892 3292
rect 16916 3290 16972 3292
rect 16996 3290 17052 3292
rect 16756 3238 16782 3290
rect 16782 3238 16812 3290
rect 16836 3238 16846 3290
rect 16846 3238 16892 3290
rect 16916 3238 16962 3290
rect 16962 3238 16972 3290
rect 16996 3238 17026 3290
rect 17026 3238 17052 3290
rect 16756 3236 16812 3238
rect 16836 3236 16892 3238
rect 16916 3236 16972 3238
rect 16996 3236 17052 3238
rect 21256 6010 21312 6012
rect 21336 6010 21392 6012
rect 21416 6010 21472 6012
rect 21496 6010 21552 6012
rect 21256 5958 21282 6010
rect 21282 5958 21312 6010
rect 21336 5958 21346 6010
rect 21346 5958 21392 6010
rect 21416 5958 21462 6010
rect 21462 5958 21472 6010
rect 21496 5958 21526 6010
rect 21526 5958 21552 6010
rect 21256 5956 21312 5958
rect 21336 5956 21392 5958
rect 21416 5956 21472 5958
rect 21496 5956 21552 5958
rect 24256 10362 24312 10364
rect 24336 10362 24392 10364
rect 24416 10362 24472 10364
rect 24496 10362 24552 10364
rect 24256 10310 24282 10362
rect 24282 10310 24312 10362
rect 24336 10310 24346 10362
rect 24346 10310 24392 10362
rect 24416 10310 24462 10362
rect 24462 10310 24472 10362
rect 24496 10310 24526 10362
rect 24526 10310 24552 10362
rect 24256 10308 24312 10310
rect 24336 10308 24392 10310
rect 24416 10308 24472 10310
rect 24496 10308 24552 10310
rect 27256 10362 27312 10364
rect 27336 10362 27392 10364
rect 27416 10362 27472 10364
rect 27496 10362 27552 10364
rect 27256 10310 27282 10362
rect 27282 10310 27312 10362
rect 27336 10310 27346 10362
rect 27346 10310 27392 10362
rect 27416 10310 27462 10362
rect 27462 10310 27472 10362
rect 27496 10310 27526 10362
rect 27526 10310 27552 10362
rect 27256 10308 27312 10310
rect 27336 10308 27392 10310
rect 27416 10308 27472 10310
rect 27496 10308 27552 10310
rect 22756 9818 22812 9820
rect 22836 9818 22892 9820
rect 22916 9818 22972 9820
rect 22996 9818 23052 9820
rect 22756 9766 22782 9818
rect 22782 9766 22812 9818
rect 22836 9766 22846 9818
rect 22846 9766 22892 9818
rect 22916 9766 22962 9818
rect 22962 9766 22972 9818
rect 22996 9766 23026 9818
rect 23026 9766 23052 9818
rect 22756 9764 22812 9766
rect 22836 9764 22892 9766
rect 22916 9764 22972 9766
rect 22996 9764 23052 9766
rect 25756 9818 25812 9820
rect 25836 9818 25892 9820
rect 25916 9818 25972 9820
rect 25996 9818 26052 9820
rect 25756 9766 25782 9818
rect 25782 9766 25812 9818
rect 25836 9766 25846 9818
rect 25846 9766 25892 9818
rect 25916 9766 25962 9818
rect 25962 9766 25972 9818
rect 25996 9766 26026 9818
rect 26026 9766 26052 9818
rect 25756 9764 25812 9766
rect 25836 9764 25892 9766
rect 25916 9764 25972 9766
rect 25996 9764 26052 9766
rect 24256 9274 24312 9276
rect 24336 9274 24392 9276
rect 24416 9274 24472 9276
rect 24496 9274 24552 9276
rect 24256 9222 24282 9274
rect 24282 9222 24312 9274
rect 24336 9222 24346 9274
rect 24346 9222 24392 9274
rect 24416 9222 24462 9274
rect 24462 9222 24472 9274
rect 24496 9222 24526 9274
rect 24526 9222 24552 9274
rect 24256 9220 24312 9222
rect 24336 9220 24392 9222
rect 24416 9220 24472 9222
rect 24496 9220 24552 9222
rect 27256 9274 27312 9276
rect 27336 9274 27392 9276
rect 27416 9274 27472 9276
rect 27496 9274 27552 9276
rect 27256 9222 27282 9274
rect 27282 9222 27312 9274
rect 27336 9222 27346 9274
rect 27346 9222 27392 9274
rect 27416 9222 27462 9274
rect 27462 9222 27472 9274
rect 27496 9222 27526 9274
rect 27526 9222 27552 9274
rect 27256 9220 27312 9222
rect 27336 9220 27392 9222
rect 27416 9220 27472 9222
rect 27496 9220 27552 9222
rect 22756 8730 22812 8732
rect 22836 8730 22892 8732
rect 22916 8730 22972 8732
rect 22996 8730 23052 8732
rect 22756 8678 22782 8730
rect 22782 8678 22812 8730
rect 22836 8678 22846 8730
rect 22846 8678 22892 8730
rect 22916 8678 22962 8730
rect 22962 8678 22972 8730
rect 22996 8678 23026 8730
rect 23026 8678 23052 8730
rect 22756 8676 22812 8678
rect 22836 8676 22892 8678
rect 22916 8676 22972 8678
rect 22996 8676 23052 8678
rect 25756 8730 25812 8732
rect 25836 8730 25892 8732
rect 25916 8730 25972 8732
rect 25996 8730 26052 8732
rect 25756 8678 25782 8730
rect 25782 8678 25812 8730
rect 25836 8678 25846 8730
rect 25846 8678 25892 8730
rect 25916 8678 25962 8730
rect 25962 8678 25972 8730
rect 25996 8678 26026 8730
rect 26026 8678 26052 8730
rect 25756 8676 25812 8678
rect 25836 8676 25892 8678
rect 25916 8676 25972 8678
rect 25996 8676 26052 8678
rect 24256 8186 24312 8188
rect 24336 8186 24392 8188
rect 24416 8186 24472 8188
rect 24496 8186 24552 8188
rect 24256 8134 24282 8186
rect 24282 8134 24312 8186
rect 24336 8134 24346 8186
rect 24346 8134 24392 8186
rect 24416 8134 24462 8186
rect 24462 8134 24472 8186
rect 24496 8134 24526 8186
rect 24526 8134 24552 8186
rect 24256 8132 24312 8134
rect 24336 8132 24392 8134
rect 24416 8132 24472 8134
rect 24496 8132 24552 8134
rect 27256 8186 27312 8188
rect 27336 8186 27392 8188
rect 27416 8186 27472 8188
rect 27496 8186 27552 8188
rect 27256 8134 27282 8186
rect 27282 8134 27312 8186
rect 27336 8134 27346 8186
rect 27346 8134 27392 8186
rect 27416 8134 27462 8186
rect 27462 8134 27472 8186
rect 27496 8134 27526 8186
rect 27526 8134 27552 8186
rect 27256 8132 27312 8134
rect 27336 8132 27392 8134
rect 27416 8132 27472 8134
rect 27496 8132 27552 8134
rect 22756 7642 22812 7644
rect 22836 7642 22892 7644
rect 22916 7642 22972 7644
rect 22996 7642 23052 7644
rect 22756 7590 22782 7642
rect 22782 7590 22812 7642
rect 22836 7590 22846 7642
rect 22846 7590 22892 7642
rect 22916 7590 22962 7642
rect 22962 7590 22972 7642
rect 22996 7590 23026 7642
rect 23026 7590 23052 7642
rect 22756 7588 22812 7590
rect 22836 7588 22892 7590
rect 22916 7588 22972 7590
rect 22996 7588 23052 7590
rect 25756 7642 25812 7644
rect 25836 7642 25892 7644
rect 25916 7642 25972 7644
rect 25996 7642 26052 7644
rect 25756 7590 25782 7642
rect 25782 7590 25812 7642
rect 25836 7590 25846 7642
rect 25846 7590 25892 7642
rect 25916 7590 25962 7642
rect 25962 7590 25972 7642
rect 25996 7590 26026 7642
rect 26026 7590 26052 7642
rect 25756 7588 25812 7590
rect 25836 7588 25892 7590
rect 25916 7588 25972 7590
rect 25996 7588 26052 7590
rect 24256 7098 24312 7100
rect 24336 7098 24392 7100
rect 24416 7098 24472 7100
rect 24496 7098 24552 7100
rect 24256 7046 24282 7098
rect 24282 7046 24312 7098
rect 24336 7046 24346 7098
rect 24346 7046 24392 7098
rect 24416 7046 24462 7098
rect 24462 7046 24472 7098
rect 24496 7046 24526 7098
rect 24526 7046 24552 7098
rect 24256 7044 24312 7046
rect 24336 7044 24392 7046
rect 24416 7044 24472 7046
rect 24496 7044 24552 7046
rect 27256 7098 27312 7100
rect 27336 7098 27392 7100
rect 27416 7098 27472 7100
rect 27496 7098 27552 7100
rect 27256 7046 27282 7098
rect 27282 7046 27312 7098
rect 27336 7046 27346 7098
rect 27346 7046 27392 7098
rect 27416 7046 27462 7098
rect 27462 7046 27472 7098
rect 27496 7046 27526 7098
rect 27526 7046 27552 7098
rect 27256 7044 27312 7046
rect 27336 7044 27392 7046
rect 27416 7044 27472 7046
rect 27496 7044 27552 7046
rect 22756 6554 22812 6556
rect 22836 6554 22892 6556
rect 22916 6554 22972 6556
rect 22996 6554 23052 6556
rect 22756 6502 22782 6554
rect 22782 6502 22812 6554
rect 22836 6502 22846 6554
rect 22846 6502 22892 6554
rect 22916 6502 22962 6554
rect 22962 6502 22972 6554
rect 22996 6502 23026 6554
rect 23026 6502 23052 6554
rect 22756 6500 22812 6502
rect 22836 6500 22892 6502
rect 22916 6500 22972 6502
rect 22996 6500 23052 6502
rect 25756 6554 25812 6556
rect 25836 6554 25892 6556
rect 25916 6554 25972 6556
rect 25996 6554 26052 6556
rect 25756 6502 25782 6554
rect 25782 6502 25812 6554
rect 25836 6502 25846 6554
rect 25846 6502 25892 6554
rect 25916 6502 25962 6554
rect 25962 6502 25972 6554
rect 25996 6502 26026 6554
rect 26026 6502 26052 6554
rect 25756 6500 25812 6502
rect 25836 6500 25892 6502
rect 25916 6500 25972 6502
rect 25996 6500 26052 6502
rect 24256 6010 24312 6012
rect 24336 6010 24392 6012
rect 24416 6010 24472 6012
rect 24496 6010 24552 6012
rect 24256 5958 24282 6010
rect 24282 5958 24312 6010
rect 24336 5958 24346 6010
rect 24346 5958 24392 6010
rect 24416 5958 24462 6010
rect 24462 5958 24472 6010
rect 24496 5958 24526 6010
rect 24526 5958 24552 6010
rect 24256 5956 24312 5958
rect 24336 5956 24392 5958
rect 24416 5956 24472 5958
rect 24496 5956 24552 5958
rect 27256 6010 27312 6012
rect 27336 6010 27392 6012
rect 27416 6010 27472 6012
rect 27496 6010 27552 6012
rect 27256 5958 27282 6010
rect 27282 5958 27312 6010
rect 27336 5958 27346 6010
rect 27346 5958 27392 6010
rect 27416 5958 27462 6010
rect 27462 5958 27472 6010
rect 27496 5958 27526 6010
rect 27526 5958 27552 6010
rect 27256 5956 27312 5958
rect 27336 5956 27392 5958
rect 27416 5956 27472 5958
rect 27496 5956 27552 5958
rect 21256 4922 21312 4924
rect 21336 4922 21392 4924
rect 21416 4922 21472 4924
rect 21496 4922 21552 4924
rect 21256 4870 21282 4922
rect 21282 4870 21312 4922
rect 21336 4870 21346 4922
rect 21346 4870 21392 4922
rect 21416 4870 21462 4922
rect 21462 4870 21472 4922
rect 21496 4870 21526 4922
rect 21526 4870 21552 4922
rect 21256 4868 21312 4870
rect 21336 4868 21392 4870
rect 21416 4868 21472 4870
rect 21496 4868 21552 4870
rect 22756 5466 22812 5468
rect 22836 5466 22892 5468
rect 22916 5466 22972 5468
rect 22996 5466 23052 5468
rect 22756 5414 22782 5466
rect 22782 5414 22812 5466
rect 22836 5414 22846 5466
rect 22846 5414 22892 5466
rect 22916 5414 22962 5466
rect 22962 5414 22972 5466
rect 22996 5414 23026 5466
rect 23026 5414 23052 5466
rect 22756 5412 22812 5414
rect 22836 5412 22892 5414
rect 22916 5412 22972 5414
rect 22996 5412 23052 5414
rect 25756 5466 25812 5468
rect 25836 5466 25892 5468
rect 25916 5466 25972 5468
rect 25996 5466 26052 5468
rect 25756 5414 25782 5466
rect 25782 5414 25812 5466
rect 25836 5414 25846 5466
rect 25846 5414 25892 5466
rect 25916 5414 25962 5466
rect 25962 5414 25972 5466
rect 25996 5414 26026 5466
rect 26026 5414 26052 5466
rect 25756 5412 25812 5414
rect 25836 5412 25892 5414
rect 25916 5412 25972 5414
rect 25996 5412 26052 5414
rect 24256 4922 24312 4924
rect 24336 4922 24392 4924
rect 24416 4922 24472 4924
rect 24496 4922 24552 4924
rect 24256 4870 24282 4922
rect 24282 4870 24312 4922
rect 24336 4870 24346 4922
rect 24346 4870 24392 4922
rect 24416 4870 24462 4922
rect 24462 4870 24472 4922
rect 24496 4870 24526 4922
rect 24526 4870 24552 4922
rect 24256 4868 24312 4870
rect 24336 4868 24392 4870
rect 24416 4868 24472 4870
rect 24496 4868 24552 4870
rect 27256 4922 27312 4924
rect 27336 4922 27392 4924
rect 27416 4922 27472 4924
rect 27496 4922 27552 4924
rect 27256 4870 27282 4922
rect 27282 4870 27312 4922
rect 27336 4870 27346 4922
rect 27346 4870 27392 4922
rect 27416 4870 27462 4922
rect 27462 4870 27472 4922
rect 27496 4870 27526 4922
rect 27526 4870 27552 4922
rect 27256 4868 27312 4870
rect 27336 4868 27392 4870
rect 27416 4868 27472 4870
rect 27496 4868 27552 4870
rect 19756 4378 19812 4380
rect 19836 4378 19892 4380
rect 19916 4378 19972 4380
rect 19996 4378 20052 4380
rect 19756 4326 19782 4378
rect 19782 4326 19812 4378
rect 19836 4326 19846 4378
rect 19846 4326 19892 4378
rect 19916 4326 19962 4378
rect 19962 4326 19972 4378
rect 19996 4326 20026 4378
rect 20026 4326 20052 4378
rect 19756 4324 19812 4326
rect 19836 4324 19892 4326
rect 19916 4324 19972 4326
rect 19996 4324 20052 4326
rect 22756 4378 22812 4380
rect 22836 4378 22892 4380
rect 22916 4378 22972 4380
rect 22996 4378 23052 4380
rect 22756 4326 22782 4378
rect 22782 4326 22812 4378
rect 22836 4326 22846 4378
rect 22846 4326 22892 4378
rect 22916 4326 22962 4378
rect 22962 4326 22972 4378
rect 22996 4326 23026 4378
rect 23026 4326 23052 4378
rect 22756 4324 22812 4326
rect 22836 4324 22892 4326
rect 22916 4324 22972 4326
rect 22996 4324 23052 4326
rect 25756 4378 25812 4380
rect 25836 4378 25892 4380
rect 25916 4378 25972 4380
rect 25996 4378 26052 4380
rect 25756 4326 25782 4378
rect 25782 4326 25812 4378
rect 25836 4326 25846 4378
rect 25846 4326 25892 4378
rect 25916 4326 25962 4378
rect 25962 4326 25972 4378
rect 25996 4326 26026 4378
rect 26026 4326 26052 4378
rect 25756 4324 25812 4326
rect 25836 4324 25892 4326
rect 25916 4324 25972 4326
rect 25996 4324 26052 4326
rect 19756 3290 19812 3292
rect 19836 3290 19892 3292
rect 19916 3290 19972 3292
rect 19996 3290 20052 3292
rect 19756 3238 19782 3290
rect 19782 3238 19812 3290
rect 19836 3238 19846 3290
rect 19846 3238 19892 3290
rect 19916 3238 19962 3290
rect 19962 3238 19972 3290
rect 19996 3238 20026 3290
rect 20026 3238 20052 3290
rect 19756 3236 19812 3238
rect 19836 3236 19892 3238
rect 19916 3236 19972 3238
rect 19996 3236 20052 3238
rect 21256 3834 21312 3836
rect 21336 3834 21392 3836
rect 21416 3834 21472 3836
rect 21496 3834 21552 3836
rect 21256 3782 21282 3834
rect 21282 3782 21312 3834
rect 21336 3782 21346 3834
rect 21346 3782 21392 3834
rect 21416 3782 21462 3834
rect 21462 3782 21472 3834
rect 21496 3782 21526 3834
rect 21526 3782 21552 3834
rect 21256 3780 21312 3782
rect 21336 3780 21392 3782
rect 21416 3780 21472 3782
rect 21496 3780 21552 3782
rect 24256 3834 24312 3836
rect 24336 3834 24392 3836
rect 24416 3834 24472 3836
rect 24496 3834 24552 3836
rect 24256 3782 24282 3834
rect 24282 3782 24312 3834
rect 24336 3782 24346 3834
rect 24346 3782 24392 3834
rect 24416 3782 24462 3834
rect 24462 3782 24472 3834
rect 24496 3782 24526 3834
rect 24526 3782 24552 3834
rect 24256 3780 24312 3782
rect 24336 3780 24392 3782
rect 24416 3780 24472 3782
rect 24496 3780 24552 3782
rect 27256 3834 27312 3836
rect 27336 3834 27392 3836
rect 27416 3834 27472 3836
rect 27496 3834 27552 3836
rect 27256 3782 27282 3834
rect 27282 3782 27312 3834
rect 27336 3782 27346 3834
rect 27346 3782 27392 3834
rect 27416 3782 27462 3834
rect 27462 3782 27472 3834
rect 27496 3782 27526 3834
rect 27526 3782 27552 3834
rect 27256 3780 27312 3782
rect 27336 3780 27392 3782
rect 27416 3780 27472 3782
rect 27496 3780 27552 3782
rect 22756 3290 22812 3292
rect 22836 3290 22892 3292
rect 22916 3290 22972 3292
rect 22996 3290 23052 3292
rect 22756 3238 22782 3290
rect 22782 3238 22812 3290
rect 22836 3238 22846 3290
rect 22846 3238 22892 3290
rect 22916 3238 22962 3290
rect 22962 3238 22972 3290
rect 22996 3238 23026 3290
rect 23026 3238 23052 3290
rect 22756 3236 22812 3238
rect 22836 3236 22892 3238
rect 22916 3236 22972 3238
rect 22996 3236 23052 3238
rect 25756 3290 25812 3292
rect 25836 3290 25892 3292
rect 25916 3290 25972 3292
rect 25996 3290 26052 3292
rect 25756 3238 25782 3290
rect 25782 3238 25812 3290
rect 25836 3238 25846 3290
rect 25846 3238 25892 3290
rect 25916 3238 25962 3290
rect 25962 3238 25972 3290
rect 25996 3238 26026 3290
rect 26026 3238 26052 3290
rect 25756 3236 25812 3238
rect 25836 3236 25892 3238
rect 25916 3236 25972 3238
rect 25996 3236 26052 3238
rect 18256 2746 18312 2748
rect 18336 2746 18392 2748
rect 18416 2746 18472 2748
rect 18496 2746 18552 2748
rect 18256 2694 18282 2746
rect 18282 2694 18312 2746
rect 18336 2694 18346 2746
rect 18346 2694 18392 2746
rect 18416 2694 18462 2746
rect 18462 2694 18472 2746
rect 18496 2694 18526 2746
rect 18526 2694 18552 2746
rect 18256 2692 18312 2694
rect 18336 2692 18392 2694
rect 18416 2692 18472 2694
rect 18496 2692 18552 2694
rect 21256 2746 21312 2748
rect 21336 2746 21392 2748
rect 21416 2746 21472 2748
rect 21496 2746 21552 2748
rect 21256 2694 21282 2746
rect 21282 2694 21312 2746
rect 21336 2694 21346 2746
rect 21346 2694 21392 2746
rect 21416 2694 21462 2746
rect 21462 2694 21472 2746
rect 21496 2694 21526 2746
rect 21526 2694 21552 2746
rect 21256 2692 21312 2694
rect 21336 2692 21392 2694
rect 21416 2692 21472 2694
rect 21496 2692 21552 2694
rect 24256 2746 24312 2748
rect 24336 2746 24392 2748
rect 24416 2746 24472 2748
rect 24496 2746 24552 2748
rect 24256 2694 24282 2746
rect 24282 2694 24312 2746
rect 24336 2694 24346 2746
rect 24346 2694 24392 2746
rect 24416 2694 24462 2746
rect 24462 2694 24472 2746
rect 24496 2694 24526 2746
rect 24526 2694 24552 2746
rect 24256 2692 24312 2694
rect 24336 2692 24392 2694
rect 24416 2692 24472 2694
rect 24496 2692 24552 2694
rect 27256 2746 27312 2748
rect 27336 2746 27392 2748
rect 27416 2746 27472 2748
rect 27496 2746 27552 2748
rect 27256 2694 27282 2746
rect 27282 2694 27312 2746
rect 27336 2694 27346 2746
rect 27346 2694 27392 2746
rect 27416 2694 27462 2746
rect 27462 2694 27472 2746
rect 27496 2694 27526 2746
rect 27526 2694 27552 2746
rect 27256 2692 27312 2694
rect 27336 2692 27392 2694
rect 27416 2692 27472 2694
rect 27496 2692 27552 2694
rect 10756 2202 10812 2204
rect 10836 2202 10892 2204
rect 10916 2202 10972 2204
rect 10996 2202 11052 2204
rect 10756 2150 10782 2202
rect 10782 2150 10812 2202
rect 10836 2150 10846 2202
rect 10846 2150 10892 2202
rect 10916 2150 10962 2202
rect 10962 2150 10972 2202
rect 10996 2150 11026 2202
rect 11026 2150 11052 2202
rect 10756 2148 10812 2150
rect 10836 2148 10892 2150
rect 10916 2148 10972 2150
rect 10996 2148 11052 2150
rect 13756 2202 13812 2204
rect 13836 2202 13892 2204
rect 13916 2202 13972 2204
rect 13996 2202 14052 2204
rect 13756 2150 13782 2202
rect 13782 2150 13812 2202
rect 13836 2150 13846 2202
rect 13846 2150 13892 2202
rect 13916 2150 13962 2202
rect 13962 2150 13972 2202
rect 13996 2150 14026 2202
rect 14026 2150 14052 2202
rect 13756 2148 13812 2150
rect 13836 2148 13892 2150
rect 13916 2148 13972 2150
rect 13996 2148 14052 2150
rect 16756 2202 16812 2204
rect 16836 2202 16892 2204
rect 16916 2202 16972 2204
rect 16996 2202 17052 2204
rect 16756 2150 16782 2202
rect 16782 2150 16812 2202
rect 16836 2150 16846 2202
rect 16846 2150 16892 2202
rect 16916 2150 16962 2202
rect 16962 2150 16972 2202
rect 16996 2150 17026 2202
rect 17026 2150 17052 2202
rect 16756 2148 16812 2150
rect 16836 2148 16892 2150
rect 16916 2148 16972 2150
rect 16996 2148 17052 2150
rect 19756 2202 19812 2204
rect 19836 2202 19892 2204
rect 19916 2202 19972 2204
rect 19996 2202 20052 2204
rect 19756 2150 19782 2202
rect 19782 2150 19812 2202
rect 19836 2150 19846 2202
rect 19846 2150 19892 2202
rect 19916 2150 19962 2202
rect 19962 2150 19972 2202
rect 19996 2150 20026 2202
rect 20026 2150 20052 2202
rect 19756 2148 19812 2150
rect 19836 2148 19892 2150
rect 19916 2148 19972 2150
rect 19996 2148 20052 2150
rect 22756 2202 22812 2204
rect 22836 2202 22892 2204
rect 22916 2202 22972 2204
rect 22996 2202 23052 2204
rect 22756 2150 22782 2202
rect 22782 2150 22812 2202
rect 22836 2150 22846 2202
rect 22846 2150 22892 2202
rect 22916 2150 22962 2202
rect 22962 2150 22972 2202
rect 22996 2150 23026 2202
rect 23026 2150 23052 2202
rect 22756 2148 22812 2150
rect 22836 2148 22892 2150
rect 22916 2148 22972 2150
rect 22996 2148 23052 2150
rect 25756 2202 25812 2204
rect 25836 2202 25892 2204
rect 25916 2202 25972 2204
rect 25996 2202 26052 2204
rect 25756 2150 25782 2202
rect 25782 2150 25812 2202
rect 25836 2150 25846 2202
rect 25846 2150 25892 2202
rect 25916 2150 25962 2202
rect 25962 2150 25972 2202
rect 25996 2150 26026 2202
rect 26026 2150 26052 2202
rect 25756 2148 25812 2150
rect 25836 2148 25892 2150
rect 25916 2148 25972 2150
rect 25996 2148 26052 2150
<< metal3 >>
rect 1744 29408 2064 29409
rect 1744 29344 1752 29408
rect 1816 29344 1832 29408
rect 1896 29344 1912 29408
rect 1976 29344 1992 29408
rect 2056 29344 2064 29408
rect 1744 29343 2064 29344
rect 4744 29408 5064 29409
rect 4744 29344 4752 29408
rect 4816 29344 4832 29408
rect 4896 29344 4912 29408
rect 4976 29344 4992 29408
rect 5056 29344 5064 29408
rect 4744 29343 5064 29344
rect 7744 29408 8064 29409
rect 7744 29344 7752 29408
rect 7816 29344 7832 29408
rect 7896 29344 7912 29408
rect 7976 29344 7992 29408
rect 8056 29344 8064 29408
rect 7744 29343 8064 29344
rect 10744 29408 11064 29409
rect 10744 29344 10752 29408
rect 10816 29344 10832 29408
rect 10896 29344 10912 29408
rect 10976 29344 10992 29408
rect 11056 29344 11064 29408
rect 10744 29343 11064 29344
rect 13744 29408 14064 29409
rect 13744 29344 13752 29408
rect 13816 29344 13832 29408
rect 13896 29344 13912 29408
rect 13976 29344 13992 29408
rect 14056 29344 14064 29408
rect 13744 29343 14064 29344
rect 16744 29408 17064 29409
rect 16744 29344 16752 29408
rect 16816 29344 16832 29408
rect 16896 29344 16912 29408
rect 16976 29344 16992 29408
rect 17056 29344 17064 29408
rect 16744 29343 17064 29344
rect 19744 29408 20064 29409
rect 19744 29344 19752 29408
rect 19816 29344 19832 29408
rect 19896 29344 19912 29408
rect 19976 29344 19992 29408
rect 20056 29344 20064 29408
rect 19744 29343 20064 29344
rect 22744 29408 23064 29409
rect 22744 29344 22752 29408
rect 22816 29344 22832 29408
rect 22896 29344 22912 29408
rect 22976 29344 22992 29408
rect 23056 29344 23064 29408
rect 22744 29343 23064 29344
rect 25744 29408 26064 29409
rect 25744 29344 25752 29408
rect 25816 29344 25832 29408
rect 25896 29344 25912 29408
rect 25976 29344 25992 29408
rect 26056 29344 26064 29408
rect 25744 29343 26064 29344
rect 3244 28864 3564 28865
rect 3244 28800 3252 28864
rect 3316 28800 3332 28864
rect 3396 28800 3412 28864
rect 3476 28800 3492 28864
rect 3556 28800 3564 28864
rect 3244 28799 3564 28800
rect 6244 28864 6564 28865
rect 6244 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6412 28864
rect 6476 28800 6492 28864
rect 6556 28800 6564 28864
rect 6244 28799 6564 28800
rect 9244 28864 9564 28865
rect 9244 28800 9252 28864
rect 9316 28800 9332 28864
rect 9396 28800 9412 28864
rect 9476 28800 9492 28864
rect 9556 28800 9564 28864
rect 9244 28799 9564 28800
rect 12244 28864 12564 28865
rect 12244 28800 12252 28864
rect 12316 28800 12332 28864
rect 12396 28800 12412 28864
rect 12476 28800 12492 28864
rect 12556 28800 12564 28864
rect 12244 28799 12564 28800
rect 15244 28864 15564 28865
rect 15244 28800 15252 28864
rect 15316 28800 15332 28864
rect 15396 28800 15412 28864
rect 15476 28800 15492 28864
rect 15556 28800 15564 28864
rect 15244 28799 15564 28800
rect 18244 28864 18564 28865
rect 18244 28800 18252 28864
rect 18316 28800 18332 28864
rect 18396 28800 18412 28864
rect 18476 28800 18492 28864
rect 18556 28800 18564 28864
rect 18244 28799 18564 28800
rect 21244 28864 21564 28865
rect 21244 28800 21252 28864
rect 21316 28800 21332 28864
rect 21396 28800 21412 28864
rect 21476 28800 21492 28864
rect 21556 28800 21564 28864
rect 21244 28799 21564 28800
rect 24244 28864 24564 28865
rect 24244 28800 24252 28864
rect 24316 28800 24332 28864
rect 24396 28800 24412 28864
rect 24476 28800 24492 28864
rect 24556 28800 24564 28864
rect 24244 28799 24564 28800
rect 27244 28864 27564 28865
rect 27244 28800 27252 28864
rect 27316 28800 27332 28864
rect 27396 28800 27412 28864
rect 27476 28800 27492 28864
rect 27556 28800 27564 28864
rect 27244 28799 27564 28800
rect 1744 28320 2064 28321
rect 1744 28256 1752 28320
rect 1816 28256 1832 28320
rect 1896 28256 1912 28320
rect 1976 28256 1992 28320
rect 2056 28256 2064 28320
rect 1744 28255 2064 28256
rect 4744 28320 5064 28321
rect 4744 28256 4752 28320
rect 4816 28256 4832 28320
rect 4896 28256 4912 28320
rect 4976 28256 4992 28320
rect 5056 28256 5064 28320
rect 4744 28255 5064 28256
rect 7744 28320 8064 28321
rect 7744 28256 7752 28320
rect 7816 28256 7832 28320
rect 7896 28256 7912 28320
rect 7976 28256 7992 28320
rect 8056 28256 8064 28320
rect 7744 28255 8064 28256
rect 10744 28320 11064 28321
rect 10744 28256 10752 28320
rect 10816 28256 10832 28320
rect 10896 28256 10912 28320
rect 10976 28256 10992 28320
rect 11056 28256 11064 28320
rect 10744 28255 11064 28256
rect 13744 28320 14064 28321
rect 13744 28256 13752 28320
rect 13816 28256 13832 28320
rect 13896 28256 13912 28320
rect 13976 28256 13992 28320
rect 14056 28256 14064 28320
rect 13744 28255 14064 28256
rect 16744 28320 17064 28321
rect 16744 28256 16752 28320
rect 16816 28256 16832 28320
rect 16896 28256 16912 28320
rect 16976 28256 16992 28320
rect 17056 28256 17064 28320
rect 16744 28255 17064 28256
rect 19744 28320 20064 28321
rect 19744 28256 19752 28320
rect 19816 28256 19832 28320
rect 19896 28256 19912 28320
rect 19976 28256 19992 28320
rect 20056 28256 20064 28320
rect 19744 28255 20064 28256
rect 22744 28320 23064 28321
rect 22744 28256 22752 28320
rect 22816 28256 22832 28320
rect 22896 28256 22912 28320
rect 22976 28256 22992 28320
rect 23056 28256 23064 28320
rect 22744 28255 23064 28256
rect 25744 28320 26064 28321
rect 25744 28256 25752 28320
rect 25816 28256 25832 28320
rect 25896 28256 25912 28320
rect 25976 28256 25992 28320
rect 26056 28256 26064 28320
rect 25744 28255 26064 28256
rect 3244 27776 3564 27777
rect 3244 27712 3252 27776
rect 3316 27712 3332 27776
rect 3396 27712 3412 27776
rect 3476 27712 3492 27776
rect 3556 27712 3564 27776
rect 3244 27711 3564 27712
rect 6244 27776 6564 27777
rect 6244 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6412 27776
rect 6476 27712 6492 27776
rect 6556 27712 6564 27776
rect 6244 27711 6564 27712
rect 9244 27776 9564 27777
rect 9244 27712 9252 27776
rect 9316 27712 9332 27776
rect 9396 27712 9412 27776
rect 9476 27712 9492 27776
rect 9556 27712 9564 27776
rect 9244 27711 9564 27712
rect 12244 27776 12564 27777
rect 12244 27712 12252 27776
rect 12316 27712 12332 27776
rect 12396 27712 12412 27776
rect 12476 27712 12492 27776
rect 12556 27712 12564 27776
rect 12244 27711 12564 27712
rect 15244 27776 15564 27777
rect 15244 27712 15252 27776
rect 15316 27712 15332 27776
rect 15396 27712 15412 27776
rect 15476 27712 15492 27776
rect 15556 27712 15564 27776
rect 15244 27711 15564 27712
rect 18244 27776 18564 27777
rect 18244 27712 18252 27776
rect 18316 27712 18332 27776
rect 18396 27712 18412 27776
rect 18476 27712 18492 27776
rect 18556 27712 18564 27776
rect 18244 27711 18564 27712
rect 21244 27776 21564 27777
rect 21244 27712 21252 27776
rect 21316 27712 21332 27776
rect 21396 27712 21412 27776
rect 21476 27712 21492 27776
rect 21556 27712 21564 27776
rect 21244 27711 21564 27712
rect 24244 27776 24564 27777
rect 24244 27712 24252 27776
rect 24316 27712 24332 27776
rect 24396 27712 24412 27776
rect 24476 27712 24492 27776
rect 24556 27712 24564 27776
rect 24244 27711 24564 27712
rect 27244 27776 27564 27777
rect 27244 27712 27252 27776
rect 27316 27712 27332 27776
rect 27396 27712 27412 27776
rect 27476 27712 27492 27776
rect 27556 27712 27564 27776
rect 27244 27711 27564 27712
rect 0 27344 800 27464
rect 1744 27232 2064 27233
rect 1744 27168 1752 27232
rect 1816 27168 1832 27232
rect 1896 27168 1912 27232
rect 1976 27168 1992 27232
rect 2056 27168 2064 27232
rect 1744 27167 2064 27168
rect 4744 27232 5064 27233
rect 4744 27168 4752 27232
rect 4816 27168 4832 27232
rect 4896 27168 4912 27232
rect 4976 27168 4992 27232
rect 5056 27168 5064 27232
rect 4744 27167 5064 27168
rect 7744 27232 8064 27233
rect 7744 27168 7752 27232
rect 7816 27168 7832 27232
rect 7896 27168 7912 27232
rect 7976 27168 7992 27232
rect 8056 27168 8064 27232
rect 7744 27167 8064 27168
rect 10744 27232 11064 27233
rect 10744 27168 10752 27232
rect 10816 27168 10832 27232
rect 10896 27168 10912 27232
rect 10976 27168 10992 27232
rect 11056 27168 11064 27232
rect 10744 27167 11064 27168
rect 13744 27232 14064 27233
rect 13744 27168 13752 27232
rect 13816 27168 13832 27232
rect 13896 27168 13912 27232
rect 13976 27168 13992 27232
rect 14056 27168 14064 27232
rect 13744 27167 14064 27168
rect 16744 27232 17064 27233
rect 16744 27168 16752 27232
rect 16816 27168 16832 27232
rect 16896 27168 16912 27232
rect 16976 27168 16992 27232
rect 17056 27168 17064 27232
rect 16744 27167 17064 27168
rect 19744 27232 20064 27233
rect 19744 27168 19752 27232
rect 19816 27168 19832 27232
rect 19896 27168 19912 27232
rect 19976 27168 19992 27232
rect 20056 27168 20064 27232
rect 19744 27167 20064 27168
rect 22744 27232 23064 27233
rect 22744 27168 22752 27232
rect 22816 27168 22832 27232
rect 22896 27168 22912 27232
rect 22976 27168 22992 27232
rect 23056 27168 23064 27232
rect 22744 27167 23064 27168
rect 25744 27232 26064 27233
rect 25744 27168 25752 27232
rect 25816 27168 25832 27232
rect 25896 27168 25912 27232
rect 25976 27168 25992 27232
rect 26056 27168 26064 27232
rect 25744 27167 26064 27168
rect 3244 26688 3564 26689
rect 3244 26624 3252 26688
rect 3316 26624 3332 26688
rect 3396 26624 3412 26688
rect 3476 26624 3492 26688
rect 3556 26624 3564 26688
rect 3244 26623 3564 26624
rect 6244 26688 6564 26689
rect 6244 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6412 26688
rect 6476 26624 6492 26688
rect 6556 26624 6564 26688
rect 6244 26623 6564 26624
rect 9244 26688 9564 26689
rect 9244 26624 9252 26688
rect 9316 26624 9332 26688
rect 9396 26624 9412 26688
rect 9476 26624 9492 26688
rect 9556 26624 9564 26688
rect 9244 26623 9564 26624
rect 12244 26688 12564 26689
rect 12244 26624 12252 26688
rect 12316 26624 12332 26688
rect 12396 26624 12412 26688
rect 12476 26624 12492 26688
rect 12556 26624 12564 26688
rect 12244 26623 12564 26624
rect 15244 26688 15564 26689
rect 15244 26624 15252 26688
rect 15316 26624 15332 26688
rect 15396 26624 15412 26688
rect 15476 26624 15492 26688
rect 15556 26624 15564 26688
rect 15244 26623 15564 26624
rect 18244 26688 18564 26689
rect 18244 26624 18252 26688
rect 18316 26624 18332 26688
rect 18396 26624 18412 26688
rect 18476 26624 18492 26688
rect 18556 26624 18564 26688
rect 18244 26623 18564 26624
rect 21244 26688 21564 26689
rect 21244 26624 21252 26688
rect 21316 26624 21332 26688
rect 21396 26624 21412 26688
rect 21476 26624 21492 26688
rect 21556 26624 21564 26688
rect 21244 26623 21564 26624
rect 24244 26688 24564 26689
rect 24244 26624 24252 26688
rect 24316 26624 24332 26688
rect 24396 26624 24412 26688
rect 24476 26624 24492 26688
rect 24556 26624 24564 26688
rect 24244 26623 24564 26624
rect 27244 26688 27564 26689
rect 27244 26624 27252 26688
rect 27316 26624 27332 26688
rect 27396 26624 27412 26688
rect 27476 26624 27492 26688
rect 27556 26624 27564 26688
rect 27244 26623 27564 26624
rect 1744 26144 2064 26145
rect 1744 26080 1752 26144
rect 1816 26080 1832 26144
rect 1896 26080 1912 26144
rect 1976 26080 1992 26144
rect 2056 26080 2064 26144
rect 1744 26079 2064 26080
rect 4744 26144 5064 26145
rect 4744 26080 4752 26144
rect 4816 26080 4832 26144
rect 4896 26080 4912 26144
rect 4976 26080 4992 26144
rect 5056 26080 5064 26144
rect 4744 26079 5064 26080
rect 7744 26144 8064 26145
rect 7744 26080 7752 26144
rect 7816 26080 7832 26144
rect 7896 26080 7912 26144
rect 7976 26080 7992 26144
rect 8056 26080 8064 26144
rect 7744 26079 8064 26080
rect 10744 26144 11064 26145
rect 10744 26080 10752 26144
rect 10816 26080 10832 26144
rect 10896 26080 10912 26144
rect 10976 26080 10992 26144
rect 11056 26080 11064 26144
rect 10744 26079 11064 26080
rect 13744 26144 14064 26145
rect 13744 26080 13752 26144
rect 13816 26080 13832 26144
rect 13896 26080 13912 26144
rect 13976 26080 13992 26144
rect 14056 26080 14064 26144
rect 13744 26079 14064 26080
rect 16744 26144 17064 26145
rect 16744 26080 16752 26144
rect 16816 26080 16832 26144
rect 16896 26080 16912 26144
rect 16976 26080 16992 26144
rect 17056 26080 17064 26144
rect 16744 26079 17064 26080
rect 19744 26144 20064 26145
rect 19744 26080 19752 26144
rect 19816 26080 19832 26144
rect 19896 26080 19912 26144
rect 19976 26080 19992 26144
rect 20056 26080 20064 26144
rect 19744 26079 20064 26080
rect 22744 26144 23064 26145
rect 22744 26080 22752 26144
rect 22816 26080 22832 26144
rect 22896 26080 22912 26144
rect 22976 26080 22992 26144
rect 23056 26080 23064 26144
rect 22744 26079 23064 26080
rect 25744 26144 26064 26145
rect 25744 26080 25752 26144
rect 25816 26080 25832 26144
rect 25896 26080 25912 26144
rect 25976 26080 25992 26144
rect 26056 26080 26064 26144
rect 25744 26079 26064 26080
rect 3244 25600 3564 25601
rect 3244 25536 3252 25600
rect 3316 25536 3332 25600
rect 3396 25536 3412 25600
rect 3476 25536 3492 25600
rect 3556 25536 3564 25600
rect 3244 25535 3564 25536
rect 6244 25600 6564 25601
rect 6244 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6412 25600
rect 6476 25536 6492 25600
rect 6556 25536 6564 25600
rect 6244 25535 6564 25536
rect 9244 25600 9564 25601
rect 9244 25536 9252 25600
rect 9316 25536 9332 25600
rect 9396 25536 9412 25600
rect 9476 25536 9492 25600
rect 9556 25536 9564 25600
rect 9244 25535 9564 25536
rect 12244 25600 12564 25601
rect 12244 25536 12252 25600
rect 12316 25536 12332 25600
rect 12396 25536 12412 25600
rect 12476 25536 12492 25600
rect 12556 25536 12564 25600
rect 12244 25535 12564 25536
rect 15244 25600 15564 25601
rect 15244 25536 15252 25600
rect 15316 25536 15332 25600
rect 15396 25536 15412 25600
rect 15476 25536 15492 25600
rect 15556 25536 15564 25600
rect 15244 25535 15564 25536
rect 18244 25600 18564 25601
rect 18244 25536 18252 25600
rect 18316 25536 18332 25600
rect 18396 25536 18412 25600
rect 18476 25536 18492 25600
rect 18556 25536 18564 25600
rect 18244 25535 18564 25536
rect 21244 25600 21564 25601
rect 21244 25536 21252 25600
rect 21316 25536 21332 25600
rect 21396 25536 21412 25600
rect 21476 25536 21492 25600
rect 21556 25536 21564 25600
rect 21244 25535 21564 25536
rect 24244 25600 24564 25601
rect 24244 25536 24252 25600
rect 24316 25536 24332 25600
rect 24396 25536 24412 25600
rect 24476 25536 24492 25600
rect 24556 25536 24564 25600
rect 24244 25535 24564 25536
rect 27244 25600 27564 25601
rect 27244 25536 27252 25600
rect 27316 25536 27332 25600
rect 27396 25536 27412 25600
rect 27476 25536 27492 25600
rect 27556 25536 27564 25600
rect 27244 25535 27564 25536
rect 1744 25056 2064 25057
rect 1744 24992 1752 25056
rect 1816 24992 1832 25056
rect 1896 24992 1912 25056
rect 1976 24992 1992 25056
rect 2056 24992 2064 25056
rect 1744 24991 2064 24992
rect 4744 25056 5064 25057
rect 4744 24992 4752 25056
rect 4816 24992 4832 25056
rect 4896 24992 4912 25056
rect 4976 24992 4992 25056
rect 5056 24992 5064 25056
rect 4744 24991 5064 24992
rect 7744 25056 8064 25057
rect 7744 24992 7752 25056
rect 7816 24992 7832 25056
rect 7896 24992 7912 25056
rect 7976 24992 7992 25056
rect 8056 24992 8064 25056
rect 7744 24991 8064 24992
rect 10744 25056 11064 25057
rect 10744 24992 10752 25056
rect 10816 24992 10832 25056
rect 10896 24992 10912 25056
rect 10976 24992 10992 25056
rect 11056 24992 11064 25056
rect 10744 24991 11064 24992
rect 13744 25056 14064 25057
rect 13744 24992 13752 25056
rect 13816 24992 13832 25056
rect 13896 24992 13912 25056
rect 13976 24992 13992 25056
rect 14056 24992 14064 25056
rect 13744 24991 14064 24992
rect 16744 25056 17064 25057
rect 16744 24992 16752 25056
rect 16816 24992 16832 25056
rect 16896 24992 16912 25056
rect 16976 24992 16992 25056
rect 17056 24992 17064 25056
rect 16744 24991 17064 24992
rect 19744 25056 20064 25057
rect 19744 24992 19752 25056
rect 19816 24992 19832 25056
rect 19896 24992 19912 25056
rect 19976 24992 19992 25056
rect 20056 24992 20064 25056
rect 19744 24991 20064 24992
rect 22744 25056 23064 25057
rect 22744 24992 22752 25056
rect 22816 24992 22832 25056
rect 22896 24992 22912 25056
rect 22976 24992 22992 25056
rect 23056 24992 23064 25056
rect 22744 24991 23064 24992
rect 25744 25056 26064 25057
rect 25744 24992 25752 25056
rect 25816 24992 25832 25056
rect 25896 24992 25912 25056
rect 25976 24992 25992 25056
rect 26056 24992 26064 25056
rect 25744 24991 26064 24992
rect 28720 24624 29520 24744
rect 3244 24512 3564 24513
rect 3244 24448 3252 24512
rect 3316 24448 3332 24512
rect 3396 24448 3412 24512
rect 3476 24448 3492 24512
rect 3556 24448 3564 24512
rect 3244 24447 3564 24448
rect 6244 24512 6564 24513
rect 6244 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6412 24512
rect 6476 24448 6492 24512
rect 6556 24448 6564 24512
rect 6244 24447 6564 24448
rect 9244 24512 9564 24513
rect 9244 24448 9252 24512
rect 9316 24448 9332 24512
rect 9396 24448 9412 24512
rect 9476 24448 9492 24512
rect 9556 24448 9564 24512
rect 9244 24447 9564 24448
rect 12244 24512 12564 24513
rect 12244 24448 12252 24512
rect 12316 24448 12332 24512
rect 12396 24448 12412 24512
rect 12476 24448 12492 24512
rect 12556 24448 12564 24512
rect 12244 24447 12564 24448
rect 15244 24512 15564 24513
rect 15244 24448 15252 24512
rect 15316 24448 15332 24512
rect 15396 24448 15412 24512
rect 15476 24448 15492 24512
rect 15556 24448 15564 24512
rect 15244 24447 15564 24448
rect 18244 24512 18564 24513
rect 18244 24448 18252 24512
rect 18316 24448 18332 24512
rect 18396 24448 18412 24512
rect 18476 24448 18492 24512
rect 18556 24448 18564 24512
rect 18244 24447 18564 24448
rect 21244 24512 21564 24513
rect 21244 24448 21252 24512
rect 21316 24448 21332 24512
rect 21396 24448 21412 24512
rect 21476 24448 21492 24512
rect 21556 24448 21564 24512
rect 21244 24447 21564 24448
rect 24244 24512 24564 24513
rect 24244 24448 24252 24512
rect 24316 24448 24332 24512
rect 24396 24448 24412 24512
rect 24476 24448 24492 24512
rect 24556 24448 24564 24512
rect 24244 24447 24564 24448
rect 27244 24512 27564 24513
rect 27244 24448 27252 24512
rect 27316 24448 27332 24512
rect 27396 24448 27412 24512
rect 27476 24448 27492 24512
rect 27556 24448 27564 24512
rect 27244 24447 27564 24448
rect 1744 23968 2064 23969
rect 1744 23904 1752 23968
rect 1816 23904 1832 23968
rect 1896 23904 1912 23968
rect 1976 23904 1992 23968
rect 2056 23904 2064 23968
rect 1744 23903 2064 23904
rect 4744 23968 5064 23969
rect 4744 23904 4752 23968
rect 4816 23904 4832 23968
rect 4896 23904 4912 23968
rect 4976 23904 4992 23968
rect 5056 23904 5064 23968
rect 4744 23903 5064 23904
rect 7744 23968 8064 23969
rect 7744 23904 7752 23968
rect 7816 23904 7832 23968
rect 7896 23904 7912 23968
rect 7976 23904 7992 23968
rect 8056 23904 8064 23968
rect 7744 23903 8064 23904
rect 10744 23968 11064 23969
rect 10744 23904 10752 23968
rect 10816 23904 10832 23968
rect 10896 23904 10912 23968
rect 10976 23904 10992 23968
rect 11056 23904 11064 23968
rect 10744 23903 11064 23904
rect 13744 23968 14064 23969
rect 13744 23904 13752 23968
rect 13816 23904 13832 23968
rect 13896 23904 13912 23968
rect 13976 23904 13992 23968
rect 14056 23904 14064 23968
rect 13744 23903 14064 23904
rect 16744 23968 17064 23969
rect 16744 23904 16752 23968
rect 16816 23904 16832 23968
rect 16896 23904 16912 23968
rect 16976 23904 16992 23968
rect 17056 23904 17064 23968
rect 16744 23903 17064 23904
rect 19744 23968 20064 23969
rect 19744 23904 19752 23968
rect 19816 23904 19832 23968
rect 19896 23904 19912 23968
rect 19976 23904 19992 23968
rect 20056 23904 20064 23968
rect 19744 23903 20064 23904
rect 22744 23968 23064 23969
rect 22744 23904 22752 23968
rect 22816 23904 22832 23968
rect 22896 23904 22912 23968
rect 22976 23904 22992 23968
rect 23056 23904 23064 23968
rect 22744 23903 23064 23904
rect 25744 23968 26064 23969
rect 25744 23904 25752 23968
rect 25816 23904 25832 23968
rect 25896 23904 25912 23968
rect 25976 23904 25992 23968
rect 26056 23904 26064 23968
rect 25744 23903 26064 23904
rect 3244 23424 3564 23425
rect 3244 23360 3252 23424
rect 3316 23360 3332 23424
rect 3396 23360 3412 23424
rect 3476 23360 3492 23424
rect 3556 23360 3564 23424
rect 3244 23359 3564 23360
rect 6244 23424 6564 23425
rect 6244 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6412 23424
rect 6476 23360 6492 23424
rect 6556 23360 6564 23424
rect 6244 23359 6564 23360
rect 9244 23424 9564 23425
rect 9244 23360 9252 23424
rect 9316 23360 9332 23424
rect 9396 23360 9412 23424
rect 9476 23360 9492 23424
rect 9556 23360 9564 23424
rect 9244 23359 9564 23360
rect 12244 23424 12564 23425
rect 12244 23360 12252 23424
rect 12316 23360 12332 23424
rect 12396 23360 12412 23424
rect 12476 23360 12492 23424
rect 12556 23360 12564 23424
rect 12244 23359 12564 23360
rect 15244 23424 15564 23425
rect 15244 23360 15252 23424
rect 15316 23360 15332 23424
rect 15396 23360 15412 23424
rect 15476 23360 15492 23424
rect 15556 23360 15564 23424
rect 15244 23359 15564 23360
rect 18244 23424 18564 23425
rect 18244 23360 18252 23424
rect 18316 23360 18332 23424
rect 18396 23360 18412 23424
rect 18476 23360 18492 23424
rect 18556 23360 18564 23424
rect 18244 23359 18564 23360
rect 21244 23424 21564 23425
rect 21244 23360 21252 23424
rect 21316 23360 21332 23424
rect 21396 23360 21412 23424
rect 21476 23360 21492 23424
rect 21556 23360 21564 23424
rect 21244 23359 21564 23360
rect 24244 23424 24564 23425
rect 24244 23360 24252 23424
rect 24316 23360 24332 23424
rect 24396 23360 24412 23424
rect 24476 23360 24492 23424
rect 24556 23360 24564 23424
rect 24244 23359 24564 23360
rect 27244 23424 27564 23425
rect 27244 23360 27252 23424
rect 27316 23360 27332 23424
rect 27396 23360 27412 23424
rect 27476 23360 27492 23424
rect 27556 23360 27564 23424
rect 27244 23359 27564 23360
rect 1744 22880 2064 22881
rect 1744 22816 1752 22880
rect 1816 22816 1832 22880
rect 1896 22816 1912 22880
rect 1976 22816 1992 22880
rect 2056 22816 2064 22880
rect 1744 22815 2064 22816
rect 4744 22880 5064 22881
rect 4744 22816 4752 22880
rect 4816 22816 4832 22880
rect 4896 22816 4912 22880
rect 4976 22816 4992 22880
rect 5056 22816 5064 22880
rect 4744 22815 5064 22816
rect 7744 22880 8064 22881
rect 7744 22816 7752 22880
rect 7816 22816 7832 22880
rect 7896 22816 7912 22880
rect 7976 22816 7992 22880
rect 8056 22816 8064 22880
rect 7744 22815 8064 22816
rect 10744 22880 11064 22881
rect 10744 22816 10752 22880
rect 10816 22816 10832 22880
rect 10896 22816 10912 22880
rect 10976 22816 10992 22880
rect 11056 22816 11064 22880
rect 10744 22815 11064 22816
rect 13744 22880 14064 22881
rect 13744 22816 13752 22880
rect 13816 22816 13832 22880
rect 13896 22816 13912 22880
rect 13976 22816 13992 22880
rect 14056 22816 14064 22880
rect 13744 22815 14064 22816
rect 16744 22880 17064 22881
rect 16744 22816 16752 22880
rect 16816 22816 16832 22880
rect 16896 22816 16912 22880
rect 16976 22816 16992 22880
rect 17056 22816 17064 22880
rect 16744 22815 17064 22816
rect 19744 22880 20064 22881
rect 19744 22816 19752 22880
rect 19816 22816 19832 22880
rect 19896 22816 19912 22880
rect 19976 22816 19992 22880
rect 20056 22816 20064 22880
rect 19744 22815 20064 22816
rect 22744 22880 23064 22881
rect 22744 22816 22752 22880
rect 22816 22816 22832 22880
rect 22896 22816 22912 22880
rect 22976 22816 22992 22880
rect 23056 22816 23064 22880
rect 22744 22815 23064 22816
rect 25744 22880 26064 22881
rect 25744 22816 25752 22880
rect 25816 22816 25832 22880
rect 25896 22816 25912 22880
rect 25976 22816 25992 22880
rect 26056 22816 26064 22880
rect 25744 22815 26064 22816
rect 3244 22336 3564 22337
rect 3244 22272 3252 22336
rect 3316 22272 3332 22336
rect 3396 22272 3412 22336
rect 3476 22272 3492 22336
rect 3556 22272 3564 22336
rect 3244 22271 3564 22272
rect 6244 22336 6564 22337
rect 6244 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6412 22336
rect 6476 22272 6492 22336
rect 6556 22272 6564 22336
rect 6244 22271 6564 22272
rect 9244 22336 9564 22337
rect 9244 22272 9252 22336
rect 9316 22272 9332 22336
rect 9396 22272 9412 22336
rect 9476 22272 9492 22336
rect 9556 22272 9564 22336
rect 9244 22271 9564 22272
rect 12244 22336 12564 22337
rect 12244 22272 12252 22336
rect 12316 22272 12332 22336
rect 12396 22272 12412 22336
rect 12476 22272 12492 22336
rect 12556 22272 12564 22336
rect 12244 22271 12564 22272
rect 15244 22336 15564 22337
rect 15244 22272 15252 22336
rect 15316 22272 15332 22336
rect 15396 22272 15412 22336
rect 15476 22272 15492 22336
rect 15556 22272 15564 22336
rect 15244 22271 15564 22272
rect 18244 22336 18564 22337
rect 18244 22272 18252 22336
rect 18316 22272 18332 22336
rect 18396 22272 18412 22336
rect 18476 22272 18492 22336
rect 18556 22272 18564 22336
rect 18244 22271 18564 22272
rect 21244 22336 21564 22337
rect 21244 22272 21252 22336
rect 21316 22272 21332 22336
rect 21396 22272 21412 22336
rect 21476 22272 21492 22336
rect 21556 22272 21564 22336
rect 21244 22271 21564 22272
rect 24244 22336 24564 22337
rect 24244 22272 24252 22336
rect 24316 22272 24332 22336
rect 24396 22272 24412 22336
rect 24476 22272 24492 22336
rect 24556 22272 24564 22336
rect 24244 22271 24564 22272
rect 27244 22336 27564 22337
rect 27244 22272 27252 22336
rect 27316 22272 27332 22336
rect 27396 22272 27412 22336
rect 27476 22272 27492 22336
rect 27556 22272 27564 22336
rect 27244 22271 27564 22272
rect 1744 21792 2064 21793
rect 1744 21728 1752 21792
rect 1816 21728 1832 21792
rect 1896 21728 1912 21792
rect 1976 21728 1992 21792
rect 2056 21728 2064 21792
rect 1744 21727 2064 21728
rect 4744 21792 5064 21793
rect 4744 21728 4752 21792
rect 4816 21728 4832 21792
rect 4896 21728 4912 21792
rect 4976 21728 4992 21792
rect 5056 21728 5064 21792
rect 4744 21727 5064 21728
rect 7744 21792 8064 21793
rect 7744 21728 7752 21792
rect 7816 21728 7832 21792
rect 7896 21728 7912 21792
rect 7976 21728 7992 21792
rect 8056 21728 8064 21792
rect 7744 21727 8064 21728
rect 10744 21792 11064 21793
rect 10744 21728 10752 21792
rect 10816 21728 10832 21792
rect 10896 21728 10912 21792
rect 10976 21728 10992 21792
rect 11056 21728 11064 21792
rect 10744 21727 11064 21728
rect 13744 21792 14064 21793
rect 13744 21728 13752 21792
rect 13816 21728 13832 21792
rect 13896 21728 13912 21792
rect 13976 21728 13992 21792
rect 14056 21728 14064 21792
rect 13744 21727 14064 21728
rect 16744 21792 17064 21793
rect 16744 21728 16752 21792
rect 16816 21728 16832 21792
rect 16896 21728 16912 21792
rect 16976 21728 16992 21792
rect 17056 21728 17064 21792
rect 16744 21727 17064 21728
rect 19744 21792 20064 21793
rect 19744 21728 19752 21792
rect 19816 21728 19832 21792
rect 19896 21728 19912 21792
rect 19976 21728 19992 21792
rect 20056 21728 20064 21792
rect 19744 21727 20064 21728
rect 22744 21792 23064 21793
rect 22744 21728 22752 21792
rect 22816 21728 22832 21792
rect 22896 21728 22912 21792
rect 22976 21728 22992 21792
rect 23056 21728 23064 21792
rect 22744 21727 23064 21728
rect 25744 21792 26064 21793
rect 25744 21728 25752 21792
rect 25816 21728 25832 21792
rect 25896 21728 25912 21792
rect 25976 21728 25992 21792
rect 26056 21728 26064 21792
rect 25744 21727 26064 21728
rect 3244 21248 3564 21249
rect 3244 21184 3252 21248
rect 3316 21184 3332 21248
rect 3396 21184 3412 21248
rect 3476 21184 3492 21248
rect 3556 21184 3564 21248
rect 3244 21183 3564 21184
rect 6244 21248 6564 21249
rect 6244 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6412 21248
rect 6476 21184 6492 21248
rect 6556 21184 6564 21248
rect 6244 21183 6564 21184
rect 9244 21248 9564 21249
rect 9244 21184 9252 21248
rect 9316 21184 9332 21248
rect 9396 21184 9412 21248
rect 9476 21184 9492 21248
rect 9556 21184 9564 21248
rect 9244 21183 9564 21184
rect 12244 21248 12564 21249
rect 12244 21184 12252 21248
rect 12316 21184 12332 21248
rect 12396 21184 12412 21248
rect 12476 21184 12492 21248
rect 12556 21184 12564 21248
rect 12244 21183 12564 21184
rect 15244 21248 15564 21249
rect 15244 21184 15252 21248
rect 15316 21184 15332 21248
rect 15396 21184 15412 21248
rect 15476 21184 15492 21248
rect 15556 21184 15564 21248
rect 15244 21183 15564 21184
rect 18244 21248 18564 21249
rect 18244 21184 18252 21248
rect 18316 21184 18332 21248
rect 18396 21184 18412 21248
rect 18476 21184 18492 21248
rect 18556 21184 18564 21248
rect 18244 21183 18564 21184
rect 21244 21248 21564 21249
rect 21244 21184 21252 21248
rect 21316 21184 21332 21248
rect 21396 21184 21412 21248
rect 21476 21184 21492 21248
rect 21556 21184 21564 21248
rect 21244 21183 21564 21184
rect 24244 21248 24564 21249
rect 24244 21184 24252 21248
rect 24316 21184 24332 21248
rect 24396 21184 24412 21248
rect 24476 21184 24492 21248
rect 24556 21184 24564 21248
rect 24244 21183 24564 21184
rect 27244 21248 27564 21249
rect 27244 21184 27252 21248
rect 27316 21184 27332 21248
rect 27396 21184 27412 21248
rect 27476 21184 27492 21248
rect 27556 21184 27564 21248
rect 27244 21183 27564 21184
rect 1744 20704 2064 20705
rect 1744 20640 1752 20704
rect 1816 20640 1832 20704
rect 1896 20640 1912 20704
rect 1976 20640 1992 20704
rect 2056 20640 2064 20704
rect 1744 20639 2064 20640
rect 4744 20704 5064 20705
rect 4744 20640 4752 20704
rect 4816 20640 4832 20704
rect 4896 20640 4912 20704
rect 4976 20640 4992 20704
rect 5056 20640 5064 20704
rect 4744 20639 5064 20640
rect 7744 20704 8064 20705
rect 7744 20640 7752 20704
rect 7816 20640 7832 20704
rect 7896 20640 7912 20704
rect 7976 20640 7992 20704
rect 8056 20640 8064 20704
rect 7744 20639 8064 20640
rect 10744 20704 11064 20705
rect 10744 20640 10752 20704
rect 10816 20640 10832 20704
rect 10896 20640 10912 20704
rect 10976 20640 10992 20704
rect 11056 20640 11064 20704
rect 10744 20639 11064 20640
rect 13744 20704 14064 20705
rect 13744 20640 13752 20704
rect 13816 20640 13832 20704
rect 13896 20640 13912 20704
rect 13976 20640 13992 20704
rect 14056 20640 14064 20704
rect 13744 20639 14064 20640
rect 16744 20704 17064 20705
rect 16744 20640 16752 20704
rect 16816 20640 16832 20704
rect 16896 20640 16912 20704
rect 16976 20640 16992 20704
rect 17056 20640 17064 20704
rect 16744 20639 17064 20640
rect 19744 20704 20064 20705
rect 19744 20640 19752 20704
rect 19816 20640 19832 20704
rect 19896 20640 19912 20704
rect 19976 20640 19992 20704
rect 20056 20640 20064 20704
rect 19744 20639 20064 20640
rect 22744 20704 23064 20705
rect 22744 20640 22752 20704
rect 22816 20640 22832 20704
rect 22896 20640 22912 20704
rect 22976 20640 22992 20704
rect 23056 20640 23064 20704
rect 22744 20639 23064 20640
rect 25744 20704 26064 20705
rect 25744 20640 25752 20704
rect 25816 20640 25832 20704
rect 25896 20640 25912 20704
rect 25976 20640 25992 20704
rect 26056 20640 26064 20704
rect 25744 20639 26064 20640
rect 3244 20160 3564 20161
rect 3244 20096 3252 20160
rect 3316 20096 3332 20160
rect 3396 20096 3412 20160
rect 3476 20096 3492 20160
rect 3556 20096 3564 20160
rect 3244 20095 3564 20096
rect 6244 20160 6564 20161
rect 6244 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6412 20160
rect 6476 20096 6492 20160
rect 6556 20096 6564 20160
rect 6244 20095 6564 20096
rect 9244 20160 9564 20161
rect 9244 20096 9252 20160
rect 9316 20096 9332 20160
rect 9396 20096 9412 20160
rect 9476 20096 9492 20160
rect 9556 20096 9564 20160
rect 9244 20095 9564 20096
rect 12244 20160 12564 20161
rect 12244 20096 12252 20160
rect 12316 20096 12332 20160
rect 12396 20096 12412 20160
rect 12476 20096 12492 20160
rect 12556 20096 12564 20160
rect 12244 20095 12564 20096
rect 15244 20160 15564 20161
rect 15244 20096 15252 20160
rect 15316 20096 15332 20160
rect 15396 20096 15412 20160
rect 15476 20096 15492 20160
rect 15556 20096 15564 20160
rect 15244 20095 15564 20096
rect 18244 20160 18564 20161
rect 18244 20096 18252 20160
rect 18316 20096 18332 20160
rect 18396 20096 18412 20160
rect 18476 20096 18492 20160
rect 18556 20096 18564 20160
rect 18244 20095 18564 20096
rect 21244 20160 21564 20161
rect 21244 20096 21252 20160
rect 21316 20096 21332 20160
rect 21396 20096 21412 20160
rect 21476 20096 21492 20160
rect 21556 20096 21564 20160
rect 21244 20095 21564 20096
rect 24244 20160 24564 20161
rect 24244 20096 24252 20160
rect 24316 20096 24332 20160
rect 24396 20096 24412 20160
rect 24476 20096 24492 20160
rect 24556 20096 24564 20160
rect 24244 20095 24564 20096
rect 27244 20160 27564 20161
rect 27244 20096 27252 20160
rect 27316 20096 27332 20160
rect 27396 20096 27412 20160
rect 27476 20096 27492 20160
rect 27556 20096 27564 20160
rect 27244 20095 27564 20096
rect 1744 19616 2064 19617
rect 1744 19552 1752 19616
rect 1816 19552 1832 19616
rect 1896 19552 1912 19616
rect 1976 19552 1992 19616
rect 2056 19552 2064 19616
rect 1744 19551 2064 19552
rect 4744 19616 5064 19617
rect 4744 19552 4752 19616
rect 4816 19552 4832 19616
rect 4896 19552 4912 19616
rect 4976 19552 4992 19616
rect 5056 19552 5064 19616
rect 4744 19551 5064 19552
rect 7744 19616 8064 19617
rect 7744 19552 7752 19616
rect 7816 19552 7832 19616
rect 7896 19552 7912 19616
rect 7976 19552 7992 19616
rect 8056 19552 8064 19616
rect 7744 19551 8064 19552
rect 10744 19616 11064 19617
rect 10744 19552 10752 19616
rect 10816 19552 10832 19616
rect 10896 19552 10912 19616
rect 10976 19552 10992 19616
rect 11056 19552 11064 19616
rect 10744 19551 11064 19552
rect 13744 19616 14064 19617
rect 13744 19552 13752 19616
rect 13816 19552 13832 19616
rect 13896 19552 13912 19616
rect 13976 19552 13992 19616
rect 14056 19552 14064 19616
rect 13744 19551 14064 19552
rect 16744 19616 17064 19617
rect 16744 19552 16752 19616
rect 16816 19552 16832 19616
rect 16896 19552 16912 19616
rect 16976 19552 16992 19616
rect 17056 19552 17064 19616
rect 16744 19551 17064 19552
rect 19744 19616 20064 19617
rect 19744 19552 19752 19616
rect 19816 19552 19832 19616
rect 19896 19552 19912 19616
rect 19976 19552 19992 19616
rect 20056 19552 20064 19616
rect 19744 19551 20064 19552
rect 22744 19616 23064 19617
rect 22744 19552 22752 19616
rect 22816 19552 22832 19616
rect 22896 19552 22912 19616
rect 22976 19552 22992 19616
rect 23056 19552 23064 19616
rect 22744 19551 23064 19552
rect 25744 19616 26064 19617
rect 25744 19552 25752 19616
rect 25816 19552 25832 19616
rect 25896 19552 25912 19616
rect 25976 19552 25992 19616
rect 26056 19552 26064 19616
rect 25744 19551 26064 19552
rect 3244 19072 3564 19073
rect 3244 19008 3252 19072
rect 3316 19008 3332 19072
rect 3396 19008 3412 19072
rect 3476 19008 3492 19072
rect 3556 19008 3564 19072
rect 3244 19007 3564 19008
rect 6244 19072 6564 19073
rect 6244 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6412 19072
rect 6476 19008 6492 19072
rect 6556 19008 6564 19072
rect 6244 19007 6564 19008
rect 9244 19072 9564 19073
rect 9244 19008 9252 19072
rect 9316 19008 9332 19072
rect 9396 19008 9412 19072
rect 9476 19008 9492 19072
rect 9556 19008 9564 19072
rect 9244 19007 9564 19008
rect 12244 19072 12564 19073
rect 12244 19008 12252 19072
rect 12316 19008 12332 19072
rect 12396 19008 12412 19072
rect 12476 19008 12492 19072
rect 12556 19008 12564 19072
rect 12244 19007 12564 19008
rect 15244 19072 15564 19073
rect 15244 19008 15252 19072
rect 15316 19008 15332 19072
rect 15396 19008 15412 19072
rect 15476 19008 15492 19072
rect 15556 19008 15564 19072
rect 15244 19007 15564 19008
rect 18244 19072 18564 19073
rect 18244 19008 18252 19072
rect 18316 19008 18332 19072
rect 18396 19008 18412 19072
rect 18476 19008 18492 19072
rect 18556 19008 18564 19072
rect 18244 19007 18564 19008
rect 21244 19072 21564 19073
rect 21244 19008 21252 19072
rect 21316 19008 21332 19072
rect 21396 19008 21412 19072
rect 21476 19008 21492 19072
rect 21556 19008 21564 19072
rect 21244 19007 21564 19008
rect 24244 19072 24564 19073
rect 24244 19008 24252 19072
rect 24316 19008 24332 19072
rect 24396 19008 24412 19072
rect 24476 19008 24492 19072
rect 24556 19008 24564 19072
rect 24244 19007 24564 19008
rect 27244 19072 27564 19073
rect 27244 19008 27252 19072
rect 27316 19008 27332 19072
rect 27396 19008 27412 19072
rect 27476 19008 27492 19072
rect 27556 19008 27564 19072
rect 27244 19007 27564 19008
rect 1744 18528 2064 18529
rect 1744 18464 1752 18528
rect 1816 18464 1832 18528
rect 1896 18464 1912 18528
rect 1976 18464 1992 18528
rect 2056 18464 2064 18528
rect 1744 18463 2064 18464
rect 4744 18528 5064 18529
rect 4744 18464 4752 18528
rect 4816 18464 4832 18528
rect 4896 18464 4912 18528
rect 4976 18464 4992 18528
rect 5056 18464 5064 18528
rect 4744 18463 5064 18464
rect 7744 18528 8064 18529
rect 7744 18464 7752 18528
rect 7816 18464 7832 18528
rect 7896 18464 7912 18528
rect 7976 18464 7992 18528
rect 8056 18464 8064 18528
rect 7744 18463 8064 18464
rect 10744 18528 11064 18529
rect 10744 18464 10752 18528
rect 10816 18464 10832 18528
rect 10896 18464 10912 18528
rect 10976 18464 10992 18528
rect 11056 18464 11064 18528
rect 10744 18463 11064 18464
rect 13744 18528 14064 18529
rect 13744 18464 13752 18528
rect 13816 18464 13832 18528
rect 13896 18464 13912 18528
rect 13976 18464 13992 18528
rect 14056 18464 14064 18528
rect 13744 18463 14064 18464
rect 16744 18528 17064 18529
rect 16744 18464 16752 18528
rect 16816 18464 16832 18528
rect 16896 18464 16912 18528
rect 16976 18464 16992 18528
rect 17056 18464 17064 18528
rect 16744 18463 17064 18464
rect 19744 18528 20064 18529
rect 19744 18464 19752 18528
rect 19816 18464 19832 18528
rect 19896 18464 19912 18528
rect 19976 18464 19992 18528
rect 20056 18464 20064 18528
rect 19744 18463 20064 18464
rect 22744 18528 23064 18529
rect 22744 18464 22752 18528
rect 22816 18464 22832 18528
rect 22896 18464 22912 18528
rect 22976 18464 22992 18528
rect 23056 18464 23064 18528
rect 22744 18463 23064 18464
rect 25744 18528 26064 18529
rect 25744 18464 25752 18528
rect 25816 18464 25832 18528
rect 25896 18464 25912 18528
rect 25976 18464 25992 18528
rect 26056 18464 26064 18528
rect 25744 18463 26064 18464
rect 3244 17984 3564 17985
rect 3244 17920 3252 17984
rect 3316 17920 3332 17984
rect 3396 17920 3412 17984
rect 3476 17920 3492 17984
rect 3556 17920 3564 17984
rect 3244 17919 3564 17920
rect 6244 17984 6564 17985
rect 6244 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6412 17984
rect 6476 17920 6492 17984
rect 6556 17920 6564 17984
rect 6244 17919 6564 17920
rect 9244 17984 9564 17985
rect 9244 17920 9252 17984
rect 9316 17920 9332 17984
rect 9396 17920 9412 17984
rect 9476 17920 9492 17984
rect 9556 17920 9564 17984
rect 9244 17919 9564 17920
rect 12244 17984 12564 17985
rect 12244 17920 12252 17984
rect 12316 17920 12332 17984
rect 12396 17920 12412 17984
rect 12476 17920 12492 17984
rect 12556 17920 12564 17984
rect 12244 17919 12564 17920
rect 15244 17984 15564 17985
rect 15244 17920 15252 17984
rect 15316 17920 15332 17984
rect 15396 17920 15412 17984
rect 15476 17920 15492 17984
rect 15556 17920 15564 17984
rect 15244 17919 15564 17920
rect 18244 17984 18564 17985
rect 18244 17920 18252 17984
rect 18316 17920 18332 17984
rect 18396 17920 18412 17984
rect 18476 17920 18492 17984
rect 18556 17920 18564 17984
rect 18244 17919 18564 17920
rect 21244 17984 21564 17985
rect 21244 17920 21252 17984
rect 21316 17920 21332 17984
rect 21396 17920 21412 17984
rect 21476 17920 21492 17984
rect 21556 17920 21564 17984
rect 21244 17919 21564 17920
rect 24244 17984 24564 17985
rect 24244 17920 24252 17984
rect 24316 17920 24332 17984
rect 24396 17920 24412 17984
rect 24476 17920 24492 17984
rect 24556 17920 24564 17984
rect 24244 17919 24564 17920
rect 27244 17984 27564 17985
rect 27244 17920 27252 17984
rect 27316 17920 27332 17984
rect 27396 17920 27412 17984
rect 27476 17920 27492 17984
rect 27556 17920 27564 17984
rect 27244 17919 27564 17920
rect 1744 17440 2064 17441
rect 1744 17376 1752 17440
rect 1816 17376 1832 17440
rect 1896 17376 1912 17440
rect 1976 17376 1992 17440
rect 2056 17376 2064 17440
rect 1744 17375 2064 17376
rect 4744 17440 5064 17441
rect 4744 17376 4752 17440
rect 4816 17376 4832 17440
rect 4896 17376 4912 17440
rect 4976 17376 4992 17440
rect 5056 17376 5064 17440
rect 4744 17375 5064 17376
rect 7744 17440 8064 17441
rect 7744 17376 7752 17440
rect 7816 17376 7832 17440
rect 7896 17376 7912 17440
rect 7976 17376 7992 17440
rect 8056 17376 8064 17440
rect 7744 17375 8064 17376
rect 10744 17440 11064 17441
rect 10744 17376 10752 17440
rect 10816 17376 10832 17440
rect 10896 17376 10912 17440
rect 10976 17376 10992 17440
rect 11056 17376 11064 17440
rect 10744 17375 11064 17376
rect 13744 17440 14064 17441
rect 13744 17376 13752 17440
rect 13816 17376 13832 17440
rect 13896 17376 13912 17440
rect 13976 17376 13992 17440
rect 14056 17376 14064 17440
rect 13744 17375 14064 17376
rect 16744 17440 17064 17441
rect 16744 17376 16752 17440
rect 16816 17376 16832 17440
rect 16896 17376 16912 17440
rect 16976 17376 16992 17440
rect 17056 17376 17064 17440
rect 16744 17375 17064 17376
rect 19744 17440 20064 17441
rect 19744 17376 19752 17440
rect 19816 17376 19832 17440
rect 19896 17376 19912 17440
rect 19976 17376 19992 17440
rect 20056 17376 20064 17440
rect 19744 17375 20064 17376
rect 22744 17440 23064 17441
rect 22744 17376 22752 17440
rect 22816 17376 22832 17440
rect 22896 17376 22912 17440
rect 22976 17376 22992 17440
rect 23056 17376 23064 17440
rect 22744 17375 23064 17376
rect 25744 17440 26064 17441
rect 25744 17376 25752 17440
rect 25816 17376 25832 17440
rect 25896 17376 25912 17440
rect 25976 17376 25992 17440
rect 26056 17376 26064 17440
rect 25744 17375 26064 17376
rect 3244 16896 3564 16897
rect 3244 16832 3252 16896
rect 3316 16832 3332 16896
rect 3396 16832 3412 16896
rect 3476 16832 3492 16896
rect 3556 16832 3564 16896
rect 3244 16831 3564 16832
rect 6244 16896 6564 16897
rect 6244 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6412 16896
rect 6476 16832 6492 16896
rect 6556 16832 6564 16896
rect 6244 16831 6564 16832
rect 9244 16896 9564 16897
rect 9244 16832 9252 16896
rect 9316 16832 9332 16896
rect 9396 16832 9412 16896
rect 9476 16832 9492 16896
rect 9556 16832 9564 16896
rect 9244 16831 9564 16832
rect 12244 16896 12564 16897
rect 12244 16832 12252 16896
rect 12316 16832 12332 16896
rect 12396 16832 12412 16896
rect 12476 16832 12492 16896
rect 12556 16832 12564 16896
rect 12244 16831 12564 16832
rect 15244 16896 15564 16897
rect 15244 16832 15252 16896
rect 15316 16832 15332 16896
rect 15396 16832 15412 16896
rect 15476 16832 15492 16896
rect 15556 16832 15564 16896
rect 15244 16831 15564 16832
rect 18244 16896 18564 16897
rect 18244 16832 18252 16896
rect 18316 16832 18332 16896
rect 18396 16832 18412 16896
rect 18476 16832 18492 16896
rect 18556 16832 18564 16896
rect 18244 16831 18564 16832
rect 21244 16896 21564 16897
rect 21244 16832 21252 16896
rect 21316 16832 21332 16896
rect 21396 16832 21412 16896
rect 21476 16832 21492 16896
rect 21556 16832 21564 16896
rect 21244 16831 21564 16832
rect 24244 16896 24564 16897
rect 24244 16832 24252 16896
rect 24316 16832 24332 16896
rect 24396 16832 24412 16896
rect 24476 16832 24492 16896
rect 24556 16832 24564 16896
rect 24244 16831 24564 16832
rect 27244 16896 27564 16897
rect 27244 16832 27252 16896
rect 27316 16832 27332 16896
rect 27396 16832 27412 16896
rect 27476 16832 27492 16896
rect 27556 16832 27564 16896
rect 27244 16831 27564 16832
rect 1744 16352 2064 16353
rect 1744 16288 1752 16352
rect 1816 16288 1832 16352
rect 1896 16288 1912 16352
rect 1976 16288 1992 16352
rect 2056 16288 2064 16352
rect 1744 16287 2064 16288
rect 4744 16352 5064 16353
rect 4744 16288 4752 16352
rect 4816 16288 4832 16352
rect 4896 16288 4912 16352
rect 4976 16288 4992 16352
rect 5056 16288 5064 16352
rect 4744 16287 5064 16288
rect 7744 16352 8064 16353
rect 7744 16288 7752 16352
rect 7816 16288 7832 16352
rect 7896 16288 7912 16352
rect 7976 16288 7992 16352
rect 8056 16288 8064 16352
rect 7744 16287 8064 16288
rect 10744 16352 11064 16353
rect 10744 16288 10752 16352
rect 10816 16288 10832 16352
rect 10896 16288 10912 16352
rect 10976 16288 10992 16352
rect 11056 16288 11064 16352
rect 10744 16287 11064 16288
rect 13744 16352 14064 16353
rect 13744 16288 13752 16352
rect 13816 16288 13832 16352
rect 13896 16288 13912 16352
rect 13976 16288 13992 16352
rect 14056 16288 14064 16352
rect 13744 16287 14064 16288
rect 16744 16352 17064 16353
rect 16744 16288 16752 16352
rect 16816 16288 16832 16352
rect 16896 16288 16912 16352
rect 16976 16288 16992 16352
rect 17056 16288 17064 16352
rect 16744 16287 17064 16288
rect 19744 16352 20064 16353
rect 19744 16288 19752 16352
rect 19816 16288 19832 16352
rect 19896 16288 19912 16352
rect 19976 16288 19992 16352
rect 20056 16288 20064 16352
rect 19744 16287 20064 16288
rect 22744 16352 23064 16353
rect 22744 16288 22752 16352
rect 22816 16288 22832 16352
rect 22896 16288 22912 16352
rect 22976 16288 22992 16352
rect 23056 16288 23064 16352
rect 22744 16287 23064 16288
rect 25744 16352 26064 16353
rect 25744 16288 25752 16352
rect 25816 16288 25832 16352
rect 25896 16288 25912 16352
rect 25976 16288 25992 16352
rect 26056 16288 26064 16352
rect 25744 16287 26064 16288
rect 3244 15808 3564 15809
rect 3244 15744 3252 15808
rect 3316 15744 3332 15808
rect 3396 15744 3412 15808
rect 3476 15744 3492 15808
rect 3556 15744 3564 15808
rect 3244 15743 3564 15744
rect 6244 15808 6564 15809
rect 6244 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6412 15808
rect 6476 15744 6492 15808
rect 6556 15744 6564 15808
rect 6244 15743 6564 15744
rect 9244 15808 9564 15809
rect 9244 15744 9252 15808
rect 9316 15744 9332 15808
rect 9396 15744 9412 15808
rect 9476 15744 9492 15808
rect 9556 15744 9564 15808
rect 9244 15743 9564 15744
rect 12244 15808 12564 15809
rect 12244 15744 12252 15808
rect 12316 15744 12332 15808
rect 12396 15744 12412 15808
rect 12476 15744 12492 15808
rect 12556 15744 12564 15808
rect 12244 15743 12564 15744
rect 15244 15808 15564 15809
rect 15244 15744 15252 15808
rect 15316 15744 15332 15808
rect 15396 15744 15412 15808
rect 15476 15744 15492 15808
rect 15556 15744 15564 15808
rect 15244 15743 15564 15744
rect 18244 15808 18564 15809
rect 18244 15744 18252 15808
rect 18316 15744 18332 15808
rect 18396 15744 18412 15808
rect 18476 15744 18492 15808
rect 18556 15744 18564 15808
rect 18244 15743 18564 15744
rect 21244 15808 21564 15809
rect 21244 15744 21252 15808
rect 21316 15744 21332 15808
rect 21396 15744 21412 15808
rect 21476 15744 21492 15808
rect 21556 15744 21564 15808
rect 21244 15743 21564 15744
rect 24244 15808 24564 15809
rect 24244 15744 24252 15808
rect 24316 15744 24332 15808
rect 24396 15744 24412 15808
rect 24476 15744 24492 15808
rect 24556 15744 24564 15808
rect 24244 15743 24564 15744
rect 27244 15808 27564 15809
rect 27244 15744 27252 15808
rect 27316 15744 27332 15808
rect 27396 15744 27412 15808
rect 27476 15744 27492 15808
rect 27556 15744 27564 15808
rect 27244 15743 27564 15744
rect 1744 15264 2064 15265
rect 1744 15200 1752 15264
rect 1816 15200 1832 15264
rect 1896 15200 1912 15264
rect 1976 15200 1992 15264
rect 2056 15200 2064 15264
rect 1744 15199 2064 15200
rect 4744 15264 5064 15265
rect 4744 15200 4752 15264
rect 4816 15200 4832 15264
rect 4896 15200 4912 15264
rect 4976 15200 4992 15264
rect 5056 15200 5064 15264
rect 4744 15199 5064 15200
rect 7744 15264 8064 15265
rect 7744 15200 7752 15264
rect 7816 15200 7832 15264
rect 7896 15200 7912 15264
rect 7976 15200 7992 15264
rect 8056 15200 8064 15264
rect 7744 15199 8064 15200
rect 10744 15264 11064 15265
rect 10744 15200 10752 15264
rect 10816 15200 10832 15264
rect 10896 15200 10912 15264
rect 10976 15200 10992 15264
rect 11056 15200 11064 15264
rect 10744 15199 11064 15200
rect 13744 15264 14064 15265
rect 13744 15200 13752 15264
rect 13816 15200 13832 15264
rect 13896 15200 13912 15264
rect 13976 15200 13992 15264
rect 14056 15200 14064 15264
rect 13744 15199 14064 15200
rect 16744 15264 17064 15265
rect 16744 15200 16752 15264
rect 16816 15200 16832 15264
rect 16896 15200 16912 15264
rect 16976 15200 16992 15264
rect 17056 15200 17064 15264
rect 16744 15199 17064 15200
rect 19744 15264 20064 15265
rect 19744 15200 19752 15264
rect 19816 15200 19832 15264
rect 19896 15200 19912 15264
rect 19976 15200 19992 15264
rect 20056 15200 20064 15264
rect 19744 15199 20064 15200
rect 22744 15264 23064 15265
rect 22744 15200 22752 15264
rect 22816 15200 22832 15264
rect 22896 15200 22912 15264
rect 22976 15200 22992 15264
rect 23056 15200 23064 15264
rect 22744 15199 23064 15200
rect 25744 15264 26064 15265
rect 25744 15200 25752 15264
rect 25816 15200 25832 15264
rect 25896 15200 25912 15264
rect 25976 15200 25992 15264
rect 26056 15200 26064 15264
rect 25744 15199 26064 15200
rect 3244 14720 3564 14721
rect 3244 14656 3252 14720
rect 3316 14656 3332 14720
rect 3396 14656 3412 14720
rect 3476 14656 3492 14720
rect 3556 14656 3564 14720
rect 3244 14655 3564 14656
rect 6244 14720 6564 14721
rect 6244 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6412 14720
rect 6476 14656 6492 14720
rect 6556 14656 6564 14720
rect 6244 14655 6564 14656
rect 9244 14720 9564 14721
rect 9244 14656 9252 14720
rect 9316 14656 9332 14720
rect 9396 14656 9412 14720
rect 9476 14656 9492 14720
rect 9556 14656 9564 14720
rect 9244 14655 9564 14656
rect 12244 14720 12564 14721
rect 12244 14656 12252 14720
rect 12316 14656 12332 14720
rect 12396 14656 12412 14720
rect 12476 14656 12492 14720
rect 12556 14656 12564 14720
rect 12244 14655 12564 14656
rect 15244 14720 15564 14721
rect 15244 14656 15252 14720
rect 15316 14656 15332 14720
rect 15396 14656 15412 14720
rect 15476 14656 15492 14720
rect 15556 14656 15564 14720
rect 15244 14655 15564 14656
rect 18244 14720 18564 14721
rect 18244 14656 18252 14720
rect 18316 14656 18332 14720
rect 18396 14656 18412 14720
rect 18476 14656 18492 14720
rect 18556 14656 18564 14720
rect 18244 14655 18564 14656
rect 21244 14720 21564 14721
rect 21244 14656 21252 14720
rect 21316 14656 21332 14720
rect 21396 14656 21412 14720
rect 21476 14656 21492 14720
rect 21556 14656 21564 14720
rect 21244 14655 21564 14656
rect 24244 14720 24564 14721
rect 24244 14656 24252 14720
rect 24316 14656 24332 14720
rect 24396 14656 24412 14720
rect 24476 14656 24492 14720
rect 24556 14656 24564 14720
rect 24244 14655 24564 14656
rect 27244 14720 27564 14721
rect 27244 14656 27252 14720
rect 27316 14656 27332 14720
rect 27396 14656 27412 14720
rect 27476 14656 27492 14720
rect 27556 14656 27564 14720
rect 27244 14655 27564 14656
rect 1744 14176 2064 14177
rect 1744 14112 1752 14176
rect 1816 14112 1832 14176
rect 1896 14112 1912 14176
rect 1976 14112 1992 14176
rect 2056 14112 2064 14176
rect 1744 14111 2064 14112
rect 4744 14176 5064 14177
rect 4744 14112 4752 14176
rect 4816 14112 4832 14176
rect 4896 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5064 14176
rect 4744 14111 5064 14112
rect 7744 14176 8064 14177
rect 7744 14112 7752 14176
rect 7816 14112 7832 14176
rect 7896 14112 7912 14176
rect 7976 14112 7992 14176
rect 8056 14112 8064 14176
rect 7744 14111 8064 14112
rect 10744 14176 11064 14177
rect 10744 14112 10752 14176
rect 10816 14112 10832 14176
rect 10896 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11064 14176
rect 10744 14111 11064 14112
rect 13744 14176 14064 14177
rect 13744 14112 13752 14176
rect 13816 14112 13832 14176
rect 13896 14112 13912 14176
rect 13976 14112 13992 14176
rect 14056 14112 14064 14176
rect 13744 14111 14064 14112
rect 16744 14176 17064 14177
rect 16744 14112 16752 14176
rect 16816 14112 16832 14176
rect 16896 14112 16912 14176
rect 16976 14112 16992 14176
rect 17056 14112 17064 14176
rect 16744 14111 17064 14112
rect 19744 14176 20064 14177
rect 19744 14112 19752 14176
rect 19816 14112 19832 14176
rect 19896 14112 19912 14176
rect 19976 14112 19992 14176
rect 20056 14112 20064 14176
rect 19744 14111 20064 14112
rect 22744 14176 23064 14177
rect 22744 14112 22752 14176
rect 22816 14112 22832 14176
rect 22896 14112 22912 14176
rect 22976 14112 22992 14176
rect 23056 14112 23064 14176
rect 22744 14111 23064 14112
rect 25744 14176 26064 14177
rect 25744 14112 25752 14176
rect 25816 14112 25832 14176
rect 25896 14112 25912 14176
rect 25976 14112 25992 14176
rect 26056 14112 26064 14176
rect 25744 14111 26064 14112
rect 0 13696 800 13728
rect 0 13640 110 13696
rect 166 13640 800 13696
rect 0 13608 800 13640
rect 3244 13632 3564 13633
rect 3244 13568 3252 13632
rect 3316 13568 3332 13632
rect 3396 13568 3412 13632
rect 3476 13568 3492 13632
rect 3556 13568 3564 13632
rect 3244 13567 3564 13568
rect 6244 13632 6564 13633
rect 6244 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6412 13632
rect 6476 13568 6492 13632
rect 6556 13568 6564 13632
rect 6244 13567 6564 13568
rect 9244 13632 9564 13633
rect 9244 13568 9252 13632
rect 9316 13568 9332 13632
rect 9396 13568 9412 13632
rect 9476 13568 9492 13632
rect 9556 13568 9564 13632
rect 9244 13567 9564 13568
rect 12244 13632 12564 13633
rect 12244 13568 12252 13632
rect 12316 13568 12332 13632
rect 12396 13568 12412 13632
rect 12476 13568 12492 13632
rect 12556 13568 12564 13632
rect 12244 13567 12564 13568
rect 15244 13632 15564 13633
rect 15244 13568 15252 13632
rect 15316 13568 15332 13632
rect 15396 13568 15412 13632
rect 15476 13568 15492 13632
rect 15556 13568 15564 13632
rect 15244 13567 15564 13568
rect 18244 13632 18564 13633
rect 18244 13568 18252 13632
rect 18316 13568 18332 13632
rect 18396 13568 18412 13632
rect 18476 13568 18492 13632
rect 18556 13568 18564 13632
rect 18244 13567 18564 13568
rect 21244 13632 21564 13633
rect 21244 13568 21252 13632
rect 21316 13568 21332 13632
rect 21396 13568 21412 13632
rect 21476 13568 21492 13632
rect 21556 13568 21564 13632
rect 21244 13567 21564 13568
rect 24244 13632 24564 13633
rect 24244 13568 24252 13632
rect 24316 13568 24332 13632
rect 24396 13568 24412 13632
rect 24476 13568 24492 13632
rect 24556 13568 24564 13632
rect 24244 13567 24564 13568
rect 27244 13632 27564 13633
rect 27244 13568 27252 13632
rect 27316 13568 27332 13632
rect 27396 13568 27412 13632
rect 27476 13568 27492 13632
rect 27556 13568 27564 13632
rect 27244 13567 27564 13568
rect 1744 13088 2064 13089
rect 1744 13024 1752 13088
rect 1816 13024 1832 13088
rect 1896 13024 1912 13088
rect 1976 13024 1992 13088
rect 2056 13024 2064 13088
rect 1744 13023 2064 13024
rect 4744 13088 5064 13089
rect 4744 13024 4752 13088
rect 4816 13024 4832 13088
rect 4896 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5064 13088
rect 4744 13023 5064 13024
rect 7744 13088 8064 13089
rect 7744 13024 7752 13088
rect 7816 13024 7832 13088
rect 7896 13024 7912 13088
rect 7976 13024 7992 13088
rect 8056 13024 8064 13088
rect 7744 13023 8064 13024
rect 10744 13088 11064 13089
rect 10744 13024 10752 13088
rect 10816 13024 10832 13088
rect 10896 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11064 13088
rect 10744 13023 11064 13024
rect 13744 13088 14064 13089
rect 13744 13024 13752 13088
rect 13816 13024 13832 13088
rect 13896 13024 13912 13088
rect 13976 13024 13992 13088
rect 14056 13024 14064 13088
rect 13744 13023 14064 13024
rect 16744 13088 17064 13089
rect 16744 13024 16752 13088
rect 16816 13024 16832 13088
rect 16896 13024 16912 13088
rect 16976 13024 16992 13088
rect 17056 13024 17064 13088
rect 16744 13023 17064 13024
rect 19744 13088 20064 13089
rect 19744 13024 19752 13088
rect 19816 13024 19832 13088
rect 19896 13024 19912 13088
rect 19976 13024 19992 13088
rect 20056 13024 20064 13088
rect 19744 13023 20064 13024
rect 22744 13088 23064 13089
rect 22744 13024 22752 13088
rect 22816 13024 22832 13088
rect 22896 13024 22912 13088
rect 22976 13024 22992 13088
rect 23056 13024 23064 13088
rect 22744 13023 23064 13024
rect 25744 13088 26064 13089
rect 25744 13024 25752 13088
rect 25816 13024 25832 13088
rect 25896 13024 25912 13088
rect 25976 13024 25992 13088
rect 26056 13024 26064 13088
rect 25744 13023 26064 13024
rect 3244 12544 3564 12545
rect 3244 12480 3252 12544
rect 3316 12480 3332 12544
rect 3396 12480 3412 12544
rect 3476 12480 3492 12544
rect 3556 12480 3564 12544
rect 3244 12479 3564 12480
rect 6244 12544 6564 12545
rect 6244 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6412 12544
rect 6476 12480 6492 12544
rect 6556 12480 6564 12544
rect 6244 12479 6564 12480
rect 9244 12544 9564 12545
rect 9244 12480 9252 12544
rect 9316 12480 9332 12544
rect 9396 12480 9412 12544
rect 9476 12480 9492 12544
rect 9556 12480 9564 12544
rect 9244 12479 9564 12480
rect 12244 12544 12564 12545
rect 12244 12480 12252 12544
rect 12316 12480 12332 12544
rect 12396 12480 12412 12544
rect 12476 12480 12492 12544
rect 12556 12480 12564 12544
rect 12244 12479 12564 12480
rect 15244 12544 15564 12545
rect 15244 12480 15252 12544
rect 15316 12480 15332 12544
rect 15396 12480 15412 12544
rect 15476 12480 15492 12544
rect 15556 12480 15564 12544
rect 15244 12479 15564 12480
rect 18244 12544 18564 12545
rect 18244 12480 18252 12544
rect 18316 12480 18332 12544
rect 18396 12480 18412 12544
rect 18476 12480 18492 12544
rect 18556 12480 18564 12544
rect 18244 12479 18564 12480
rect 21244 12544 21564 12545
rect 21244 12480 21252 12544
rect 21316 12480 21332 12544
rect 21396 12480 21412 12544
rect 21476 12480 21492 12544
rect 21556 12480 21564 12544
rect 21244 12479 21564 12480
rect 24244 12544 24564 12545
rect 24244 12480 24252 12544
rect 24316 12480 24332 12544
rect 24396 12480 24412 12544
rect 24476 12480 24492 12544
rect 24556 12480 24564 12544
rect 24244 12479 24564 12480
rect 27244 12544 27564 12545
rect 27244 12480 27252 12544
rect 27316 12480 27332 12544
rect 27396 12480 27412 12544
rect 27476 12480 27492 12544
rect 27556 12480 27564 12544
rect 27244 12479 27564 12480
rect 105 12202 171 12205
rect 23473 12202 23539 12205
rect 105 12200 23539 12202
rect 105 12144 110 12200
rect 166 12144 23478 12200
rect 23534 12144 23539 12200
rect 105 12142 23539 12144
rect 105 12139 171 12142
rect 23473 12139 23539 12142
rect 1744 12000 2064 12001
rect 1744 11936 1752 12000
rect 1816 11936 1832 12000
rect 1896 11936 1912 12000
rect 1976 11936 1992 12000
rect 2056 11936 2064 12000
rect 1744 11935 2064 11936
rect 4744 12000 5064 12001
rect 4744 11936 4752 12000
rect 4816 11936 4832 12000
rect 4896 11936 4912 12000
rect 4976 11936 4992 12000
rect 5056 11936 5064 12000
rect 4744 11935 5064 11936
rect 7744 12000 8064 12001
rect 7744 11936 7752 12000
rect 7816 11936 7832 12000
rect 7896 11936 7912 12000
rect 7976 11936 7992 12000
rect 8056 11936 8064 12000
rect 7744 11935 8064 11936
rect 10744 12000 11064 12001
rect 10744 11936 10752 12000
rect 10816 11936 10832 12000
rect 10896 11936 10912 12000
rect 10976 11936 10992 12000
rect 11056 11936 11064 12000
rect 10744 11935 11064 11936
rect 13744 12000 14064 12001
rect 13744 11936 13752 12000
rect 13816 11936 13832 12000
rect 13896 11936 13912 12000
rect 13976 11936 13992 12000
rect 14056 11936 14064 12000
rect 13744 11935 14064 11936
rect 16744 12000 17064 12001
rect 16744 11936 16752 12000
rect 16816 11936 16832 12000
rect 16896 11936 16912 12000
rect 16976 11936 16992 12000
rect 17056 11936 17064 12000
rect 16744 11935 17064 11936
rect 19744 12000 20064 12001
rect 19744 11936 19752 12000
rect 19816 11936 19832 12000
rect 19896 11936 19912 12000
rect 19976 11936 19992 12000
rect 20056 11936 20064 12000
rect 19744 11935 20064 11936
rect 22744 12000 23064 12001
rect 22744 11936 22752 12000
rect 22816 11936 22832 12000
rect 22896 11936 22912 12000
rect 22976 11936 22992 12000
rect 23056 11936 23064 12000
rect 22744 11935 23064 11936
rect 25744 12000 26064 12001
rect 25744 11936 25752 12000
rect 25816 11936 25832 12000
rect 25896 11936 25912 12000
rect 25976 11936 25992 12000
rect 26056 11936 26064 12000
rect 25744 11935 26064 11936
rect 18413 11794 18479 11797
rect 19333 11794 19399 11797
rect 18413 11792 19399 11794
rect 18413 11736 18418 11792
rect 18474 11736 19338 11792
rect 19394 11736 19399 11792
rect 18413 11734 19399 11736
rect 18413 11731 18479 11734
rect 19333 11731 19399 11734
rect 3244 11456 3564 11457
rect 3244 11392 3252 11456
rect 3316 11392 3332 11456
rect 3396 11392 3412 11456
rect 3476 11392 3492 11456
rect 3556 11392 3564 11456
rect 3244 11391 3564 11392
rect 6244 11456 6564 11457
rect 6244 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6412 11456
rect 6476 11392 6492 11456
rect 6556 11392 6564 11456
rect 6244 11391 6564 11392
rect 9244 11456 9564 11457
rect 9244 11392 9252 11456
rect 9316 11392 9332 11456
rect 9396 11392 9412 11456
rect 9476 11392 9492 11456
rect 9556 11392 9564 11456
rect 9244 11391 9564 11392
rect 12244 11456 12564 11457
rect 12244 11392 12252 11456
rect 12316 11392 12332 11456
rect 12396 11392 12412 11456
rect 12476 11392 12492 11456
rect 12556 11392 12564 11456
rect 12244 11391 12564 11392
rect 15244 11456 15564 11457
rect 15244 11392 15252 11456
rect 15316 11392 15332 11456
rect 15396 11392 15412 11456
rect 15476 11392 15492 11456
rect 15556 11392 15564 11456
rect 15244 11391 15564 11392
rect 18244 11456 18564 11457
rect 18244 11392 18252 11456
rect 18316 11392 18332 11456
rect 18396 11392 18412 11456
rect 18476 11392 18492 11456
rect 18556 11392 18564 11456
rect 18244 11391 18564 11392
rect 21244 11456 21564 11457
rect 21244 11392 21252 11456
rect 21316 11392 21332 11456
rect 21396 11392 21412 11456
rect 21476 11392 21492 11456
rect 21556 11392 21564 11456
rect 21244 11391 21564 11392
rect 24244 11456 24564 11457
rect 24244 11392 24252 11456
rect 24316 11392 24332 11456
rect 24396 11392 24412 11456
rect 24476 11392 24492 11456
rect 24556 11392 24564 11456
rect 24244 11391 24564 11392
rect 27244 11456 27564 11457
rect 27244 11392 27252 11456
rect 27316 11392 27332 11456
rect 27396 11392 27412 11456
rect 27476 11392 27492 11456
rect 27556 11392 27564 11456
rect 27244 11391 27564 11392
rect 28720 11117 29520 11144
rect 28717 11114 29520 11117
rect 28636 11112 29520 11114
rect 28636 11056 28722 11112
rect 28778 11056 29520 11112
rect 28636 11054 29520 11056
rect 28717 11051 29520 11054
rect 28720 11024 29520 11051
rect 1744 10912 2064 10913
rect 1744 10848 1752 10912
rect 1816 10848 1832 10912
rect 1896 10848 1912 10912
rect 1976 10848 1992 10912
rect 2056 10848 2064 10912
rect 1744 10847 2064 10848
rect 4744 10912 5064 10913
rect 4744 10848 4752 10912
rect 4816 10848 4832 10912
rect 4896 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5064 10912
rect 4744 10847 5064 10848
rect 7744 10912 8064 10913
rect 7744 10848 7752 10912
rect 7816 10848 7832 10912
rect 7896 10848 7912 10912
rect 7976 10848 7992 10912
rect 8056 10848 8064 10912
rect 7744 10847 8064 10848
rect 10744 10912 11064 10913
rect 10744 10848 10752 10912
rect 10816 10848 10832 10912
rect 10896 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11064 10912
rect 10744 10847 11064 10848
rect 13744 10912 14064 10913
rect 13744 10848 13752 10912
rect 13816 10848 13832 10912
rect 13896 10848 13912 10912
rect 13976 10848 13992 10912
rect 14056 10848 14064 10912
rect 13744 10847 14064 10848
rect 16744 10912 17064 10913
rect 16744 10848 16752 10912
rect 16816 10848 16832 10912
rect 16896 10848 16912 10912
rect 16976 10848 16992 10912
rect 17056 10848 17064 10912
rect 16744 10847 17064 10848
rect 19744 10912 20064 10913
rect 19744 10848 19752 10912
rect 19816 10848 19832 10912
rect 19896 10848 19912 10912
rect 19976 10848 19992 10912
rect 20056 10848 20064 10912
rect 19744 10847 20064 10848
rect 22744 10912 23064 10913
rect 22744 10848 22752 10912
rect 22816 10848 22832 10912
rect 22896 10848 22912 10912
rect 22976 10848 22992 10912
rect 23056 10848 23064 10912
rect 22744 10847 23064 10848
rect 25744 10912 26064 10913
rect 25744 10848 25752 10912
rect 25816 10848 25832 10912
rect 25896 10848 25912 10912
rect 25976 10848 25992 10912
rect 26056 10848 26064 10912
rect 25744 10847 26064 10848
rect 3244 10368 3564 10369
rect 3244 10304 3252 10368
rect 3316 10304 3332 10368
rect 3396 10304 3412 10368
rect 3476 10304 3492 10368
rect 3556 10304 3564 10368
rect 3244 10303 3564 10304
rect 6244 10368 6564 10369
rect 6244 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6412 10368
rect 6476 10304 6492 10368
rect 6556 10304 6564 10368
rect 6244 10303 6564 10304
rect 9244 10368 9564 10369
rect 9244 10304 9252 10368
rect 9316 10304 9332 10368
rect 9396 10304 9412 10368
rect 9476 10304 9492 10368
rect 9556 10304 9564 10368
rect 9244 10303 9564 10304
rect 12244 10368 12564 10369
rect 12244 10304 12252 10368
rect 12316 10304 12332 10368
rect 12396 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12564 10368
rect 12244 10303 12564 10304
rect 15244 10368 15564 10369
rect 15244 10304 15252 10368
rect 15316 10304 15332 10368
rect 15396 10304 15412 10368
rect 15476 10304 15492 10368
rect 15556 10304 15564 10368
rect 15244 10303 15564 10304
rect 18244 10368 18564 10369
rect 18244 10304 18252 10368
rect 18316 10304 18332 10368
rect 18396 10304 18412 10368
rect 18476 10304 18492 10368
rect 18556 10304 18564 10368
rect 18244 10303 18564 10304
rect 21244 10368 21564 10369
rect 21244 10304 21252 10368
rect 21316 10304 21332 10368
rect 21396 10304 21412 10368
rect 21476 10304 21492 10368
rect 21556 10304 21564 10368
rect 21244 10303 21564 10304
rect 24244 10368 24564 10369
rect 24244 10304 24252 10368
rect 24316 10304 24332 10368
rect 24396 10304 24412 10368
rect 24476 10304 24492 10368
rect 24556 10304 24564 10368
rect 24244 10303 24564 10304
rect 27244 10368 27564 10369
rect 27244 10304 27252 10368
rect 27316 10304 27332 10368
rect 27396 10304 27412 10368
rect 27476 10304 27492 10368
rect 27556 10304 27564 10368
rect 27244 10303 27564 10304
rect 1744 9824 2064 9825
rect 1744 9760 1752 9824
rect 1816 9760 1832 9824
rect 1896 9760 1912 9824
rect 1976 9760 1992 9824
rect 2056 9760 2064 9824
rect 1744 9759 2064 9760
rect 4744 9824 5064 9825
rect 4744 9760 4752 9824
rect 4816 9760 4832 9824
rect 4896 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5064 9824
rect 4744 9759 5064 9760
rect 7744 9824 8064 9825
rect 7744 9760 7752 9824
rect 7816 9760 7832 9824
rect 7896 9760 7912 9824
rect 7976 9760 7992 9824
rect 8056 9760 8064 9824
rect 7744 9759 8064 9760
rect 10744 9824 11064 9825
rect 10744 9760 10752 9824
rect 10816 9760 10832 9824
rect 10896 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11064 9824
rect 10744 9759 11064 9760
rect 13744 9824 14064 9825
rect 13744 9760 13752 9824
rect 13816 9760 13832 9824
rect 13896 9760 13912 9824
rect 13976 9760 13992 9824
rect 14056 9760 14064 9824
rect 13744 9759 14064 9760
rect 16744 9824 17064 9825
rect 16744 9760 16752 9824
rect 16816 9760 16832 9824
rect 16896 9760 16912 9824
rect 16976 9760 16992 9824
rect 17056 9760 17064 9824
rect 16744 9759 17064 9760
rect 19744 9824 20064 9825
rect 19744 9760 19752 9824
rect 19816 9760 19832 9824
rect 19896 9760 19912 9824
rect 19976 9760 19992 9824
rect 20056 9760 20064 9824
rect 19744 9759 20064 9760
rect 22744 9824 23064 9825
rect 22744 9760 22752 9824
rect 22816 9760 22832 9824
rect 22896 9760 22912 9824
rect 22976 9760 22992 9824
rect 23056 9760 23064 9824
rect 22744 9759 23064 9760
rect 25744 9824 26064 9825
rect 25744 9760 25752 9824
rect 25816 9760 25832 9824
rect 25896 9760 25912 9824
rect 25976 9760 25992 9824
rect 26056 9760 26064 9824
rect 25744 9759 26064 9760
rect 3244 9280 3564 9281
rect 3244 9216 3252 9280
rect 3316 9216 3332 9280
rect 3396 9216 3412 9280
rect 3476 9216 3492 9280
rect 3556 9216 3564 9280
rect 3244 9215 3564 9216
rect 6244 9280 6564 9281
rect 6244 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6412 9280
rect 6476 9216 6492 9280
rect 6556 9216 6564 9280
rect 6244 9215 6564 9216
rect 9244 9280 9564 9281
rect 9244 9216 9252 9280
rect 9316 9216 9332 9280
rect 9396 9216 9412 9280
rect 9476 9216 9492 9280
rect 9556 9216 9564 9280
rect 9244 9215 9564 9216
rect 12244 9280 12564 9281
rect 12244 9216 12252 9280
rect 12316 9216 12332 9280
rect 12396 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12564 9280
rect 12244 9215 12564 9216
rect 15244 9280 15564 9281
rect 15244 9216 15252 9280
rect 15316 9216 15332 9280
rect 15396 9216 15412 9280
rect 15476 9216 15492 9280
rect 15556 9216 15564 9280
rect 15244 9215 15564 9216
rect 18244 9280 18564 9281
rect 18244 9216 18252 9280
rect 18316 9216 18332 9280
rect 18396 9216 18412 9280
rect 18476 9216 18492 9280
rect 18556 9216 18564 9280
rect 18244 9215 18564 9216
rect 21244 9280 21564 9281
rect 21244 9216 21252 9280
rect 21316 9216 21332 9280
rect 21396 9216 21412 9280
rect 21476 9216 21492 9280
rect 21556 9216 21564 9280
rect 21244 9215 21564 9216
rect 24244 9280 24564 9281
rect 24244 9216 24252 9280
rect 24316 9216 24332 9280
rect 24396 9216 24412 9280
rect 24476 9216 24492 9280
rect 24556 9216 24564 9280
rect 24244 9215 24564 9216
rect 27244 9280 27564 9281
rect 27244 9216 27252 9280
rect 27316 9216 27332 9280
rect 27396 9216 27412 9280
rect 27476 9216 27492 9280
rect 27556 9216 27564 9280
rect 27244 9215 27564 9216
rect 1744 8736 2064 8737
rect 1744 8672 1752 8736
rect 1816 8672 1832 8736
rect 1896 8672 1912 8736
rect 1976 8672 1992 8736
rect 2056 8672 2064 8736
rect 1744 8671 2064 8672
rect 4744 8736 5064 8737
rect 4744 8672 4752 8736
rect 4816 8672 4832 8736
rect 4896 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5064 8736
rect 4744 8671 5064 8672
rect 7744 8736 8064 8737
rect 7744 8672 7752 8736
rect 7816 8672 7832 8736
rect 7896 8672 7912 8736
rect 7976 8672 7992 8736
rect 8056 8672 8064 8736
rect 7744 8671 8064 8672
rect 10744 8736 11064 8737
rect 10744 8672 10752 8736
rect 10816 8672 10832 8736
rect 10896 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11064 8736
rect 10744 8671 11064 8672
rect 13744 8736 14064 8737
rect 13744 8672 13752 8736
rect 13816 8672 13832 8736
rect 13896 8672 13912 8736
rect 13976 8672 13992 8736
rect 14056 8672 14064 8736
rect 13744 8671 14064 8672
rect 16744 8736 17064 8737
rect 16744 8672 16752 8736
rect 16816 8672 16832 8736
rect 16896 8672 16912 8736
rect 16976 8672 16992 8736
rect 17056 8672 17064 8736
rect 16744 8671 17064 8672
rect 19744 8736 20064 8737
rect 19744 8672 19752 8736
rect 19816 8672 19832 8736
rect 19896 8672 19912 8736
rect 19976 8672 19992 8736
rect 20056 8672 20064 8736
rect 19744 8671 20064 8672
rect 22744 8736 23064 8737
rect 22744 8672 22752 8736
rect 22816 8672 22832 8736
rect 22896 8672 22912 8736
rect 22976 8672 22992 8736
rect 23056 8672 23064 8736
rect 22744 8671 23064 8672
rect 25744 8736 26064 8737
rect 25744 8672 25752 8736
rect 25816 8672 25832 8736
rect 25896 8672 25912 8736
rect 25976 8672 25992 8736
rect 26056 8672 26064 8736
rect 25744 8671 26064 8672
rect 3244 8192 3564 8193
rect 3244 8128 3252 8192
rect 3316 8128 3332 8192
rect 3396 8128 3412 8192
rect 3476 8128 3492 8192
rect 3556 8128 3564 8192
rect 3244 8127 3564 8128
rect 6244 8192 6564 8193
rect 6244 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6412 8192
rect 6476 8128 6492 8192
rect 6556 8128 6564 8192
rect 6244 8127 6564 8128
rect 9244 8192 9564 8193
rect 9244 8128 9252 8192
rect 9316 8128 9332 8192
rect 9396 8128 9412 8192
rect 9476 8128 9492 8192
rect 9556 8128 9564 8192
rect 9244 8127 9564 8128
rect 12244 8192 12564 8193
rect 12244 8128 12252 8192
rect 12316 8128 12332 8192
rect 12396 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12564 8192
rect 12244 8127 12564 8128
rect 15244 8192 15564 8193
rect 15244 8128 15252 8192
rect 15316 8128 15332 8192
rect 15396 8128 15412 8192
rect 15476 8128 15492 8192
rect 15556 8128 15564 8192
rect 15244 8127 15564 8128
rect 18244 8192 18564 8193
rect 18244 8128 18252 8192
rect 18316 8128 18332 8192
rect 18396 8128 18412 8192
rect 18476 8128 18492 8192
rect 18556 8128 18564 8192
rect 18244 8127 18564 8128
rect 21244 8192 21564 8193
rect 21244 8128 21252 8192
rect 21316 8128 21332 8192
rect 21396 8128 21412 8192
rect 21476 8128 21492 8192
rect 21556 8128 21564 8192
rect 21244 8127 21564 8128
rect 24244 8192 24564 8193
rect 24244 8128 24252 8192
rect 24316 8128 24332 8192
rect 24396 8128 24412 8192
rect 24476 8128 24492 8192
rect 24556 8128 24564 8192
rect 24244 8127 24564 8128
rect 27244 8192 27564 8193
rect 27244 8128 27252 8192
rect 27316 8128 27332 8192
rect 27396 8128 27412 8192
rect 27476 8128 27492 8192
rect 27556 8128 27564 8192
rect 27244 8127 27564 8128
rect 1744 7648 2064 7649
rect 1744 7584 1752 7648
rect 1816 7584 1832 7648
rect 1896 7584 1912 7648
rect 1976 7584 1992 7648
rect 2056 7584 2064 7648
rect 1744 7583 2064 7584
rect 4744 7648 5064 7649
rect 4744 7584 4752 7648
rect 4816 7584 4832 7648
rect 4896 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5064 7648
rect 4744 7583 5064 7584
rect 7744 7648 8064 7649
rect 7744 7584 7752 7648
rect 7816 7584 7832 7648
rect 7896 7584 7912 7648
rect 7976 7584 7992 7648
rect 8056 7584 8064 7648
rect 7744 7583 8064 7584
rect 10744 7648 11064 7649
rect 10744 7584 10752 7648
rect 10816 7584 10832 7648
rect 10896 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11064 7648
rect 10744 7583 11064 7584
rect 13744 7648 14064 7649
rect 13744 7584 13752 7648
rect 13816 7584 13832 7648
rect 13896 7584 13912 7648
rect 13976 7584 13992 7648
rect 14056 7584 14064 7648
rect 13744 7583 14064 7584
rect 16744 7648 17064 7649
rect 16744 7584 16752 7648
rect 16816 7584 16832 7648
rect 16896 7584 16912 7648
rect 16976 7584 16992 7648
rect 17056 7584 17064 7648
rect 16744 7583 17064 7584
rect 19744 7648 20064 7649
rect 19744 7584 19752 7648
rect 19816 7584 19832 7648
rect 19896 7584 19912 7648
rect 19976 7584 19992 7648
rect 20056 7584 20064 7648
rect 19744 7583 20064 7584
rect 22744 7648 23064 7649
rect 22744 7584 22752 7648
rect 22816 7584 22832 7648
rect 22896 7584 22912 7648
rect 22976 7584 22992 7648
rect 23056 7584 23064 7648
rect 22744 7583 23064 7584
rect 25744 7648 26064 7649
rect 25744 7584 25752 7648
rect 25816 7584 25832 7648
rect 25896 7584 25912 7648
rect 25976 7584 25992 7648
rect 26056 7584 26064 7648
rect 25744 7583 26064 7584
rect 3244 7104 3564 7105
rect 3244 7040 3252 7104
rect 3316 7040 3332 7104
rect 3396 7040 3412 7104
rect 3476 7040 3492 7104
rect 3556 7040 3564 7104
rect 3244 7039 3564 7040
rect 6244 7104 6564 7105
rect 6244 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6412 7104
rect 6476 7040 6492 7104
rect 6556 7040 6564 7104
rect 6244 7039 6564 7040
rect 9244 7104 9564 7105
rect 9244 7040 9252 7104
rect 9316 7040 9332 7104
rect 9396 7040 9412 7104
rect 9476 7040 9492 7104
rect 9556 7040 9564 7104
rect 9244 7039 9564 7040
rect 12244 7104 12564 7105
rect 12244 7040 12252 7104
rect 12316 7040 12332 7104
rect 12396 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12564 7104
rect 12244 7039 12564 7040
rect 15244 7104 15564 7105
rect 15244 7040 15252 7104
rect 15316 7040 15332 7104
rect 15396 7040 15412 7104
rect 15476 7040 15492 7104
rect 15556 7040 15564 7104
rect 15244 7039 15564 7040
rect 18244 7104 18564 7105
rect 18244 7040 18252 7104
rect 18316 7040 18332 7104
rect 18396 7040 18412 7104
rect 18476 7040 18492 7104
rect 18556 7040 18564 7104
rect 18244 7039 18564 7040
rect 21244 7104 21564 7105
rect 21244 7040 21252 7104
rect 21316 7040 21332 7104
rect 21396 7040 21412 7104
rect 21476 7040 21492 7104
rect 21556 7040 21564 7104
rect 21244 7039 21564 7040
rect 24244 7104 24564 7105
rect 24244 7040 24252 7104
rect 24316 7040 24332 7104
rect 24396 7040 24412 7104
rect 24476 7040 24492 7104
rect 24556 7040 24564 7104
rect 24244 7039 24564 7040
rect 27244 7104 27564 7105
rect 27244 7040 27252 7104
rect 27316 7040 27332 7104
rect 27396 7040 27412 7104
rect 27476 7040 27492 7104
rect 27556 7040 27564 7104
rect 27244 7039 27564 7040
rect 1744 6560 2064 6561
rect 1744 6496 1752 6560
rect 1816 6496 1832 6560
rect 1896 6496 1912 6560
rect 1976 6496 1992 6560
rect 2056 6496 2064 6560
rect 1744 6495 2064 6496
rect 4744 6560 5064 6561
rect 4744 6496 4752 6560
rect 4816 6496 4832 6560
rect 4896 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5064 6560
rect 4744 6495 5064 6496
rect 7744 6560 8064 6561
rect 7744 6496 7752 6560
rect 7816 6496 7832 6560
rect 7896 6496 7912 6560
rect 7976 6496 7992 6560
rect 8056 6496 8064 6560
rect 7744 6495 8064 6496
rect 10744 6560 11064 6561
rect 10744 6496 10752 6560
rect 10816 6496 10832 6560
rect 10896 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11064 6560
rect 10744 6495 11064 6496
rect 13744 6560 14064 6561
rect 13744 6496 13752 6560
rect 13816 6496 13832 6560
rect 13896 6496 13912 6560
rect 13976 6496 13992 6560
rect 14056 6496 14064 6560
rect 13744 6495 14064 6496
rect 16744 6560 17064 6561
rect 16744 6496 16752 6560
rect 16816 6496 16832 6560
rect 16896 6496 16912 6560
rect 16976 6496 16992 6560
rect 17056 6496 17064 6560
rect 16744 6495 17064 6496
rect 19744 6560 20064 6561
rect 19744 6496 19752 6560
rect 19816 6496 19832 6560
rect 19896 6496 19912 6560
rect 19976 6496 19992 6560
rect 20056 6496 20064 6560
rect 19744 6495 20064 6496
rect 22744 6560 23064 6561
rect 22744 6496 22752 6560
rect 22816 6496 22832 6560
rect 22896 6496 22912 6560
rect 22976 6496 22992 6560
rect 23056 6496 23064 6560
rect 22744 6495 23064 6496
rect 25744 6560 26064 6561
rect 25744 6496 25752 6560
rect 25816 6496 25832 6560
rect 25896 6496 25912 6560
rect 25976 6496 25992 6560
rect 26056 6496 26064 6560
rect 25744 6495 26064 6496
rect 3244 6016 3564 6017
rect 3244 5952 3252 6016
rect 3316 5952 3332 6016
rect 3396 5952 3412 6016
rect 3476 5952 3492 6016
rect 3556 5952 3564 6016
rect 3244 5951 3564 5952
rect 6244 6016 6564 6017
rect 6244 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6412 6016
rect 6476 5952 6492 6016
rect 6556 5952 6564 6016
rect 6244 5951 6564 5952
rect 9244 6016 9564 6017
rect 9244 5952 9252 6016
rect 9316 5952 9332 6016
rect 9396 5952 9412 6016
rect 9476 5952 9492 6016
rect 9556 5952 9564 6016
rect 9244 5951 9564 5952
rect 12244 6016 12564 6017
rect 12244 5952 12252 6016
rect 12316 5952 12332 6016
rect 12396 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12564 6016
rect 12244 5951 12564 5952
rect 15244 6016 15564 6017
rect 15244 5952 15252 6016
rect 15316 5952 15332 6016
rect 15396 5952 15412 6016
rect 15476 5952 15492 6016
rect 15556 5952 15564 6016
rect 15244 5951 15564 5952
rect 18244 6016 18564 6017
rect 18244 5952 18252 6016
rect 18316 5952 18332 6016
rect 18396 5952 18412 6016
rect 18476 5952 18492 6016
rect 18556 5952 18564 6016
rect 18244 5951 18564 5952
rect 21244 6016 21564 6017
rect 21244 5952 21252 6016
rect 21316 5952 21332 6016
rect 21396 5952 21412 6016
rect 21476 5952 21492 6016
rect 21556 5952 21564 6016
rect 21244 5951 21564 5952
rect 24244 6016 24564 6017
rect 24244 5952 24252 6016
rect 24316 5952 24332 6016
rect 24396 5952 24412 6016
rect 24476 5952 24492 6016
rect 24556 5952 24564 6016
rect 24244 5951 24564 5952
rect 27244 6016 27564 6017
rect 27244 5952 27252 6016
rect 27316 5952 27332 6016
rect 27396 5952 27412 6016
rect 27476 5952 27492 6016
rect 27556 5952 27564 6016
rect 27244 5951 27564 5952
rect 1744 5472 2064 5473
rect 1744 5408 1752 5472
rect 1816 5408 1832 5472
rect 1896 5408 1912 5472
rect 1976 5408 1992 5472
rect 2056 5408 2064 5472
rect 1744 5407 2064 5408
rect 4744 5472 5064 5473
rect 4744 5408 4752 5472
rect 4816 5408 4832 5472
rect 4896 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5064 5472
rect 4744 5407 5064 5408
rect 7744 5472 8064 5473
rect 7744 5408 7752 5472
rect 7816 5408 7832 5472
rect 7896 5408 7912 5472
rect 7976 5408 7992 5472
rect 8056 5408 8064 5472
rect 7744 5407 8064 5408
rect 10744 5472 11064 5473
rect 10744 5408 10752 5472
rect 10816 5408 10832 5472
rect 10896 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11064 5472
rect 10744 5407 11064 5408
rect 13744 5472 14064 5473
rect 13744 5408 13752 5472
rect 13816 5408 13832 5472
rect 13896 5408 13912 5472
rect 13976 5408 13992 5472
rect 14056 5408 14064 5472
rect 13744 5407 14064 5408
rect 16744 5472 17064 5473
rect 16744 5408 16752 5472
rect 16816 5408 16832 5472
rect 16896 5408 16912 5472
rect 16976 5408 16992 5472
rect 17056 5408 17064 5472
rect 16744 5407 17064 5408
rect 19744 5472 20064 5473
rect 19744 5408 19752 5472
rect 19816 5408 19832 5472
rect 19896 5408 19912 5472
rect 19976 5408 19992 5472
rect 20056 5408 20064 5472
rect 19744 5407 20064 5408
rect 22744 5472 23064 5473
rect 22744 5408 22752 5472
rect 22816 5408 22832 5472
rect 22896 5408 22912 5472
rect 22976 5408 22992 5472
rect 23056 5408 23064 5472
rect 22744 5407 23064 5408
rect 25744 5472 26064 5473
rect 25744 5408 25752 5472
rect 25816 5408 25832 5472
rect 25896 5408 25912 5472
rect 25976 5408 25992 5472
rect 26056 5408 26064 5472
rect 25744 5407 26064 5408
rect 3244 4928 3564 4929
rect 3244 4864 3252 4928
rect 3316 4864 3332 4928
rect 3396 4864 3412 4928
rect 3476 4864 3492 4928
rect 3556 4864 3564 4928
rect 3244 4863 3564 4864
rect 6244 4928 6564 4929
rect 6244 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6412 4928
rect 6476 4864 6492 4928
rect 6556 4864 6564 4928
rect 6244 4863 6564 4864
rect 9244 4928 9564 4929
rect 9244 4864 9252 4928
rect 9316 4864 9332 4928
rect 9396 4864 9412 4928
rect 9476 4864 9492 4928
rect 9556 4864 9564 4928
rect 9244 4863 9564 4864
rect 12244 4928 12564 4929
rect 12244 4864 12252 4928
rect 12316 4864 12332 4928
rect 12396 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12564 4928
rect 12244 4863 12564 4864
rect 15244 4928 15564 4929
rect 15244 4864 15252 4928
rect 15316 4864 15332 4928
rect 15396 4864 15412 4928
rect 15476 4864 15492 4928
rect 15556 4864 15564 4928
rect 15244 4863 15564 4864
rect 18244 4928 18564 4929
rect 18244 4864 18252 4928
rect 18316 4864 18332 4928
rect 18396 4864 18412 4928
rect 18476 4864 18492 4928
rect 18556 4864 18564 4928
rect 18244 4863 18564 4864
rect 21244 4928 21564 4929
rect 21244 4864 21252 4928
rect 21316 4864 21332 4928
rect 21396 4864 21412 4928
rect 21476 4864 21492 4928
rect 21556 4864 21564 4928
rect 21244 4863 21564 4864
rect 24244 4928 24564 4929
rect 24244 4864 24252 4928
rect 24316 4864 24332 4928
rect 24396 4864 24412 4928
rect 24476 4864 24492 4928
rect 24556 4864 24564 4928
rect 24244 4863 24564 4864
rect 27244 4928 27564 4929
rect 27244 4864 27252 4928
rect 27316 4864 27332 4928
rect 27396 4864 27412 4928
rect 27476 4864 27492 4928
rect 27556 4864 27564 4928
rect 27244 4863 27564 4864
rect 1744 4384 2064 4385
rect 1744 4320 1752 4384
rect 1816 4320 1832 4384
rect 1896 4320 1912 4384
rect 1976 4320 1992 4384
rect 2056 4320 2064 4384
rect 1744 4319 2064 4320
rect 4744 4384 5064 4385
rect 4744 4320 4752 4384
rect 4816 4320 4832 4384
rect 4896 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5064 4384
rect 4744 4319 5064 4320
rect 7744 4384 8064 4385
rect 7744 4320 7752 4384
rect 7816 4320 7832 4384
rect 7896 4320 7912 4384
rect 7976 4320 7992 4384
rect 8056 4320 8064 4384
rect 7744 4319 8064 4320
rect 10744 4384 11064 4385
rect 10744 4320 10752 4384
rect 10816 4320 10832 4384
rect 10896 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11064 4384
rect 10744 4319 11064 4320
rect 13744 4384 14064 4385
rect 13744 4320 13752 4384
rect 13816 4320 13832 4384
rect 13896 4320 13912 4384
rect 13976 4320 13992 4384
rect 14056 4320 14064 4384
rect 13744 4319 14064 4320
rect 16744 4384 17064 4385
rect 16744 4320 16752 4384
rect 16816 4320 16832 4384
rect 16896 4320 16912 4384
rect 16976 4320 16992 4384
rect 17056 4320 17064 4384
rect 16744 4319 17064 4320
rect 19744 4384 20064 4385
rect 19744 4320 19752 4384
rect 19816 4320 19832 4384
rect 19896 4320 19912 4384
rect 19976 4320 19992 4384
rect 20056 4320 20064 4384
rect 19744 4319 20064 4320
rect 22744 4384 23064 4385
rect 22744 4320 22752 4384
rect 22816 4320 22832 4384
rect 22896 4320 22912 4384
rect 22976 4320 22992 4384
rect 23056 4320 23064 4384
rect 22744 4319 23064 4320
rect 25744 4384 26064 4385
rect 25744 4320 25752 4384
rect 25816 4320 25832 4384
rect 25896 4320 25912 4384
rect 25976 4320 25992 4384
rect 26056 4320 26064 4384
rect 25744 4319 26064 4320
rect 7649 4042 7715 4045
rect 10041 4042 10107 4045
rect 7649 4040 10107 4042
rect 7649 3984 7654 4040
rect 7710 3984 10046 4040
rect 10102 3984 10107 4040
rect 7649 3982 10107 3984
rect 7649 3979 7715 3982
rect 10041 3979 10107 3982
rect 3244 3840 3564 3841
rect 3244 3776 3252 3840
rect 3316 3776 3332 3840
rect 3396 3776 3412 3840
rect 3476 3776 3492 3840
rect 3556 3776 3564 3840
rect 3244 3775 3564 3776
rect 6244 3840 6564 3841
rect 6244 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6412 3840
rect 6476 3776 6492 3840
rect 6556 3776 6564 3840
rect 6244 3775 6564 3776
rect 9244 3840 9564 3841
rect 9244 3776 9252 3840
rect 9316 3776 9332 3840
rect 9396 3776 9412 3840
rect 9476 3776 9492 3840
rect 9556 3776 9564 3840
rect 9244 3775 9564 3776
rect 12244 3840 12564 3841
rect 12244 3776 12252 3840
rect 12316 3776 12332 3840
rect 12396 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12564 3840
rect 12244 3775 12564 3776
rect 15244 3840 15564 3841
rect 15244 3776 15252 3840
rect 15316 3776 15332 3840
rect 15396 3776 15412 3840
rect 15476 3776 15492 3840
rect 15556 3776 15564 3840
rect 15244 3775 15564 3776
rect 18244 3840 18564 3841
rect 18244 3776 18252 3840
rect 18316 3776 18332 3840
rect 18396 3776 18412 3840
rect 18476 3776 18492 3840
rect 18556 3776 18564 3840
rect 18244 3775 18564 3776
rect 21244 3840 21564 3841
rect 21244 3776 21252 3840
rect 21316 3776 21332 3840
rect 21396 3776 21412 3840
rect 21476 3776 21492 3840
rect 21556 3776 21564 3840
rect 21244 3775 21564 3776
rect 24244 3840 24564 3841
rect 24244 3776 24252 3840
rect 24316 3776 24332 3840
rect 24396 3776 24412 3840
rect 24476 3776 24492 3840
rect 24556 3776 24564 3840
rect 24244 3775 24564 3776
rect 27244 3840 27564 3841
rect 27244 3776 27252 3840
rect 27316 3776 27332 3840
rect 27396 3776 27412 3840
rect 27476 3776 27492 3840
rect 27556 3776 27564 3840
rect 27244 3775 27564 3776
rect 1744 3296 2064 3297
rect 1744 3232 1752 3296
rect 1816 3232 1832 3296
rect 1896 3232 1912 3296
rect 1976 3232 1992 3296
rect 2056 3232 2064 3296
rect 1744 3231 2064 3232
rect 4744 3296 5064 3297
rect 4744 3232 4752 3296
rect 4816 3232 4832 3296
rect 4896 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5064 3296
rect 4744 3231 5064 3232
rect 7744 3296 8064 3297
rect 7744 3232 7752 3296
rect 7816 3232 7832 3296
rect 7896 3232 7912 3296
rect 7976 3232 7992 3296
rect 8056 3232 8064 3296
rect 7744 3231 8064 3232
rect 10744 3296 11064 3297
rect 10744 3232 10752 3296
rect 10816 3232 10832 3296
rect 10896 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11064 3296
rect 10744 3231 11064 3232
rect 13744 3296 14064 3297
rect 13744 3232 13752 3296
rect 13816 3232 13832 3296
rect 13896 3232 13912 3296
rect 13976 3232 13992 3296
rect 14056 3232 14064 3296
rect 13744 3231 14064 3232
rect 16744 3296 17064 3297
rect 16744 3232 16752 3296
rect 16816 3232 16832 3296
rect 16896 3232 16912 3296
rect 16976 3232 16992 3296
rect 17056 3232 17064 3296
rect 16744 3231 17064 3232
rect 19744 3296 20064 3297
rect 19744 3232 19752 3296
rect 19816 3232 19832 3296
rect 19896 3232 19912 3296
rect 19976 3232 19992 3296
rect 20056 3232 20064 3296
rect 19744 3231 20064 3232
rect 22744 3296 23064 3297
rect 22744 3232 22752 3296
rect 22816 3232 22832 3296
rect 22896 3232 22912 3296
rect 22976 3232 22992 3296
rect 23056 3232 23064 3296
rect 22744 3231 23064 3232
rect 25744 3296 26064 3297
rect 25744 3232 25752 3296
rect 25816 3232 25832 3296
rect 25896 3232 25912 3296
rect 25976 3232 25992 3296
rect 26056 3232 26064 3296
rect 25744 3231 26064 3232
rect 3244 2752 3564 2753
rect 3244 2688 3252 2752
rect 3316 2688 3332 2752
rect 3396 2688 3412 2752
rect 3476 2688 3492 2752
rect 3556 2688 3564 2752
rect 3244 2687 3564 2688
rect 6244 2752 6564 2753
rect 6244 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6412 2752
rect 6476 2688 6492 2752
rect 6556 2688 6564 2752
rect 6244 2687 6564 2688
rect 9244 2752 9564 2753
rect 9244 2688 9252 2752
rect 9316 2688 9332 2752
rect 9396 2688 9412 2752
rect 9476 2688 9492 2752
rect 9556 2688 9564 2752
rect 9244 2687 9564 2688
rect 12244 2752 12564 2753
rect 12244 2688 12252 2752
rect 12316 2688 12332 2752
rect 12396 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12564 2752
rect 12244 2687 12564 2688
rect 15244 2752 15564 2753
rect 15244 2688 15252 2752
rect 15316 2688 15332 2752
rect 15396 2688 15412 2752
rect 15476 2688 15492 2752
rect 15556 2688 15564 2752
rect 15244 2687 15564 2688
rect 18244 2752 18564 2753
rect 18244 2688 18252 2752
rect 18316 2688 18332 2752
rect 18396 2688 18412 2752
rect 18476 2688 18492 2752
rect 18556 2688 18564 2752
rect 18244 2687 18564 2688
rect 21244 2752 21564 2753
rect 21244 2688 21252 2752
rect 21316 2688 21332 2752
rect 21396 2688 21412 2752
rect 21476 2688 21492 2752
rect 21556 2688 21564 2752
rect 21244 2687 21564 2688
rect 24244 2752 24564 2753
rect 24244 2688 24252 2752
rect 24316 2688 24332 2752
rect 24396 2688 24412 2752
rect 24476 2688 24492 2752
rect 24556 2688 24564 2752
rect 24244 2687 24564 2688
rect 27244 2752 27564 2753
rect 27244 2688 27252 2752
rect 27316 2688 27332 2752
rect 27396 2688 27412 2752
rect 27476 2688 27492 2752
rect 27556 2688 27564 2752
rect 27244 2687 27564 2688
rect 10041 2546 10107 2549
rect 14365 2546 14431 2549
rect 10041 2544 14431 2546
rect 10041 2488 10046 2544
rect 10102 2488 14370 2544
rect 14426 2488 14431 2544
rect 10041 2486 14431 2488
rect 10041 2483 10107 2486
rect 14365 2483 14431 2486
rect 1744 2208 2064 2209
rect 1744 2144 1752 2208
rect 1816 2144 1832 2208
rect 1896 2144 1912 2208
rect 1976 2144 1992 2208
rect 2056 2144 2064 2208
rect 1744 2143 2064 2144
rect 4744 2208 5064 2209
rect 4744 2144 4752 2208
rect 4816 2144 4832 2208
rect 4896 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5064 2208
rect 4744 2143 5064 2144
rect 7744 2208 8064 2209
rect 7744 2144 7752 2208
rect 7816 2144 7832 2208
rect 7896 2144 7912 2208
rect 7976 2144 7992 2208
rect 8056 2144 8064 2208
rect 7744 2143 8064 2144
rect 10744 2208 11064 2209
rect 10744 2144 10752 2208
rect 10816 2144 10832 2208
rect 10896 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11064 2208
rect 10744 2143 11064 2144
rect 13744 2208 14064 2209
rect 13744 2144 13752 2208
rect 13816 2144 13832 2208
rect 13896 2144 13912 2208
rect 13976 2144 13992 2208
rect 14056 2144 14064 2208
rect 13744 2143 14064 2144
rect 16744 2208 17064 2209
rect 16744 2144 16752 2208
rect 16816 2144 16832 2208
rect 16896 2144 16912 2208
rect 16976 2144 16992 2208
rect 17056 2144 17064 2208
rect 16744 2143 17064 2144
rect 19744 2208 20064 2209
rect 19744 2144 19752 2208
rect 19816 2144 19832 2208
rect 19896 2144 19912 2208
rect 19976 2144 19992 2208
rect 20056 2144 20064 2208
rect 19744 2143 20064 2144
rect 22744 2208 23064 2209
rect 22744 2144 22752 2208
rect 22816 2144 22832 2208
rect 22896 2144 22912 2208
rect 22976 2144 22992 2208
rect 23056 2144 23064 2208
rect 22744 2143 23064 2144
rect 25744 2208 26064 2209
rect 25744 2144 25752 2208
rect 25816 2144 25832 2208
rect 25896 2144 25912 2208
rect 25976 2144 25992 2208
rect 26056 2144 26064 2208
rect 25744 2143 26064 2144
<< via3 >>
rect 1752 29404 1816 29408
rect 1752 29348 1756 29404
rect 1756 29348 1812 29404
rect 1812 29348 1816 29404
rect 1752 29344 1816 29348
rect 1832 29404 1896 29408
rect 1832 29348 1836 29404
rect 1836 29348 1892 29404
rect 1892 29348 1896 29404
rect 1832 29344 1896 29348
rect 1912 29404 1976 29408
rect 1912 29348 1916 29404
rect 1916 29348 1972 29404
rect 1972 29348 1976 29404
rect 1912 29344 1976 29348
rect 1992 29404 2056 29408
rect 1992 29348 1996 29404
rect 1996 29348 2052 29404
rect 2052 29348 2056 29404
rect 1992 29344 2056 29348
rect 4752 29404 4816 29408
rect 4752 29348 4756 29404
rect 4756 29348 4812 29404
rect 4812 29348 4816 29404
rect 4752 29344 4816 29348
rect 4832 29404 4896 29408
rect 4832 29348 4836 29404
rect 4836 29348 4892 29404
rect 4892 29348 4896 29404
rect 4832 29344 4896 29348
rect 4912 29404 4976 29408
rect 4912 29348 4916 29404
rect 4916 29348 4972 29404
rect 4972 29348 4976 29404
rect 4912 29344 4976 29348
rect 4992 29404 5056 29408
rect 4992 29348 4996 29404
rect 4996 29348 5052 29404
rect 5052 29348 5056 29404
rect 4992 29344 5056 29348
rect 7752 29404 7816 29408
rect 7752 29348 7756 29404
rect 7756 29348 7812 29404
rect 7812 29348 7816 29404
rect 7752 29344 7816 29348
rect 7832 29404 7896 29408
rect 7832 29348 7836 29404
rect 7836 29348 7892 29404
rect 7892 29348 7896 29404
rect 7832 29344 7896 29348
rect 7912 29404 7976 29408
rect 7912 29348 7916 29404
rect 7916 29348 7972 29404
rect 7972 29348 7976 29404
rect 7912 29344 7976 29348
rect 7992 29404 8056 29408
rect 7992 29348 7996 29404
rect 7996 29348 8052 29404
rect 8052 29348 8056 29404
rect 7992 29344 8056 29348
rect 10752 29404 10816 29408
rect 10752 29348 10756 29404
rect 10756 29348 10812 29404
rect 10812 29348 10816 29404
rect 10752 29344 10816 29348
rect 10832 29404 10896 29408
rect 10832 29348 10836 29404
rect 10836 29348 10892 29404
rect 10892 29348 10896 29404
rect 10832 29344 10896 29348
rect 10912 29404 10976 29408
rect 10912 29348 10916 29404
rect 10916 29348 10972 29404
rect 10972 29348 10976 29404
rect 10912 29344 10976 29348
rect 10992 29404 11056 29408
rect 10992 29348 10996 29404
rect 10996 29348 11052 29404
rect 11052 29348 11056 29404
rect 10992 29344 11056 29348
rect 13752 29404 13816 29408
rect 13752 29348 13756 29404
rect 13756 29348 13812 29404
rect 13812 29348 13816 29404
rect 13752 29344 13816 29348
rect 13832 29404 13896 29408
rect 13832 29348 13836 29404
rect 13836 29348 13892 29404
rect 13892 29348 13896 29404
rect 13832 29344 13896 29348
rect 13912 29404 13976 29408
rect 13912 29348 13916 29404
rect 13916 29348 13972 29404
rect 13972 29348 13976 29404
rect 13912 29344 13976 29348
rect 13992 29404 14056 29408
rect 13992 29348 13996 29404
rect 13996 29348 14052 29404
rect 14052 29348 14056 29404
rect 13992 29344 14056 29348
rect 16752 29404 16816 29408
rect 16752 29348 16756 29404
rect 16756 29348 16812 29404
rect 16812 29348 16816 29404
rect 16752 29344 16816 29348
rect 16832 29404 16896 29408
rect 16832 29348 16836 29404
rect 16836 29348 16892 29404
rect 16892 29348 16896 29404
rect 16832 29344 16896 29348
rect 16912 29404 16976 29408
rect 16912 29348 16916 29404
rect 16916 29348 16972 29404
rect 16972 29348 16976 29404
rect 16912 29344 16976 29348
rect 16992 29404 17056 29408
rect 16992 29348 16996 29404
rect 16996 29348 17052 29404
rect 17052 29348 17056 29404
rect 16992 29344 17056 29348
rect 19752 29404 19816 29408
rect 19752 29348 19756 29404
rect 19756 29348 19812 29404
rect 19812 29348 19816 29404
rect 19752 29344 19816 29348
rect 19832 29404 19896 29408
rect 19832 29348 19836 29404
rect 19836 29348 19892 29404
rect 19892 29348 19896 29404
rect 19832 29344 19896 29348
rect 19912 29404 19976 29408
rect 19912 29348 19916 29404
rect 19916 29348 19972 29404
rect 19972 29348 19976 29404
rect 19912 29344 19976 29348
rect 19992 29404 20056 29408
rect 19992 29348 19996 29404
rect 19996 29348 20052 29404
rect 20052 29348 20056 29404
rect 19992 29344 20056 29348
rect 22752 29404 22816 29408
rect 22752 29348 22756 29404
rect 22756 29348 22812 29404
rect 22812 29348 22816 29404
rect 22752 29344 22816 29348
rect 22832 29404 22896 29408
rect 22832 29348 22836 29404
rect 22836 29348 22892 29404
rect 22892 29348 22896 29404
rect 22832 29344 22896 29348
rect 22912 29404 22976 29408
rect 22912 29348 22916 29404
rect 22916 29348 22972 29404
rect 22972 29348 22976 29404
rect 22912 29344 22976 29348
rect 22992 29404 23056 29408
rect 22992 29348 22996 29404
rect 22996 29348 23052 29404
rect 23052 29348 23056 29404
rect 22992 29344 23056 29348
rect 25752 29404 25816 29408
rect 25752 29348 25756 29404
rect 25756 29348 25812 29404
rect 25812 29348 25816 29404
rect 25752 29344 25816 29348
rect 25832 29404 25896 29408
rect 25832 29348 25836 29404
rect 25836 29348 25892 29404
rect 25892 29348 25896 29404
rect 25832 29344 25896 29348
rect 25912 29404 25976 29408
rect 25912 29348 25916 29404
rect 25916 29348 25972 29404
rect 25972 29348 25976 29404
rect 25912 29344 25976 29348
rect 25992 29404 26056 29408
rect 25992 29348 25996 29404
rect 25996 29348 26052 29404
rect 26052 29348 26056 29404
rect 25992 29344 26056 29348
rect 3252 28860 3316 28864
rect 3252 28804 3256 28860
rect 3256 28804 3312 28860
rect 3312 28804 3316 28860
rect 3252 28800 3316 28804
rect 3332 28860 3396 28864
rect 3332 28804 3336 28860
rect 3336 28804 3392 28860
rect 3392 28804 3396 28860
rect 3332 28800 3396 28804
rect 3412 28860 3476 28864
rect 3412 28804 3416 28860
rect 3416 28804 3472 28860
rect 3472 28804 3476 28860
rect 3412 28800 3476 28804
rect 3492 28860 3556 28864
rect 3492 28804 3496 28860
rect 3496 28804 3552 28860
rect 3552 28804 3556 28860
rect 3492 28800 3556 28804
rect 6252 28860 6316 28864
rect 6252 28804 6256 28860
rect 6256 28804 6312 28860
rect 6312 28804 6316 28860
rect 6252 28800 6316 28804
rect 6332 28860 6396 28864
rect 6332 28804 6336 28860
rect 6336 28804 6392 28860
rect 6392 28804 6396 28860
rect 6332 28800 6396 28804
rect 6412 28860 6476 28864
rect 6412 28804 6416 28860
rect 6416 28804 6472 28860
rect 6472 28804 6476 28860
rect 6412 28800 6476 28804
rect 6492 28860 6556 28864
rect 6492 28804 6496 28860
rect 6496 28804 6552 28860
rect 6552 28804 6556 28860
rect 6492 28800 6556 28804
rect 9252 28860 9316 28864
rect 9252 28804 9256 28860
rect 9256 28804 9312 28860
rect 9312 28804 9316 28860
rect 9252 28800 9316 28804
rect 9332 28860 9396 28864
rect 9332 28804 9336 28860
rect 9336 28804 9392 28860
rect 9392 28804 9396 28860
rect 9332 28800 9396 28804
rect 9412 28860 9476 28864
rect 9412 28804 9416 28860
rect 9416 28804 9472 28860
rect 9472 28804 9476 28860
rect 9412 28800 9476 28804
rect 9492 28860 9556 28864
rect 9492 28804 9496 28860
rect 9496 28804 9552 28860
rect 9552 28804 9556 28860
rect 9492 28800 9556 28804
rect 12252 28860 12316 28864
rect 12252 28804 12256 28860
rect 12256 28804 12312 28860
rect 12312 28804 12316 28860
rect 12252 28800 12316 28804
rect 12332 28860 12396 28864
rect 12332 28804 12336 28860
rect 12336 28804 12392 28860
rect 12392 28804 12396 28860
rect 12332 28800 12396 28804
rect 12412 28860 12476 28864
rect 12412 28804 12416 28860
rect 12416 28804 12472 28860
rect 12472 28804 12476 28860
rect 12412 28800 12476 28804
rect 12492 28860 12556 28864
rect 12492 28804 12496 28860
rect 12496 28804 12552 28860
rect 12552 28804 12556 28860
rect 12492 28800 12556 28804
rect 15252 28860 15316 28864
rect 15252 28804 15256 28860
rect 15256 28804 15312 28860
rect 15312 28804 15316 28860
rect 15252 28800 15316 28804
rect 15332 28860 15396 28864
rect 15332 28804 15336 28860
rect 15336 28804 15392 28860
rect 15392 28804 15396 28860
rect 15332 28800 15396 28804
rect 15412 28860 15476 28864
rect 15412 28804 15416 28860
rect 15416 28804 15472 28860
rect 15472 28804 15476 28860
rect 15412 28800 15476 28804
rect 15492 28860 15556 28864
rect 15492 28804 15496 28860
rect 15496 28804 15552 28860
rect 15552 28804 15556 28860
rect 15492 28800 15556 28804
rect 18252 28860 18316 28864
rect 18252 28804 18256 28860
rect 18256 28804 18312 28860
rect 18312 28804 18316 28860
rect 18252 28800 18316 28804
rect 18332 28860 18396 28864
rect 18332 28804 18336 28860
rect 18336 28804 18392 28860
rect 18392 28804 18396 28860
rect 18332 28800 18396 28804
rect 18412 28860 18476 28864
rect 18412 28804 18416 28860
rect 18416 28804 18472 28860
rect 18472 28804 18476 28860
rect 18412 28800 18476 28804
rect 18492 28860 18556 28864
rect 18492 28804 18496 28860
rect 18496 28804 18552 28860
rect 18552 28804 18556 28860
rect 18492 28800 18556 28804
rect 21252 28860 21316 28864
rect 21252 28804 21256 28860
rect 21256 28804 21312 28860
rect 21312 28804 21316 28860
rect 21252 28800 21316 28804
rect 21332 28860 21396 28864
rect 21332 28804 21336 28860
rect 21336 28804 21392 28860
rect 21392 28804 21396 28860
rect 21332 28800 21396 28804
rect 21412 28860 21476 28864
rect 21412 28804 21416 28860
rect 21416 28804 21472 28860
rect 21472 28804 21476 28860
rect 21412 28800 21476 28804
rect 21492 28860 21556 28864
rect 21492 28804 21496 28860
rect 21496 28804 21552 28860
rect 21552 28804 21556 28860
rect 21492 28800 21556 28804
rect 24252 28860 24316 28864
rect 24252 28804 24256 28860
rect 24256 28804 24312 28860
rect 24312 28804 24316 28860
rect 24252 28800 24316 28804
rect 24332 28860 24396 28864
rect 24332 28804 24336 28860
rect 24336 28804 24392 28860
rect 24392 28804 24396 28860
rect 24332 28800 24396 28804
rect 24412 28860 24476 28864
rect 24412 28804 24416 28860
rect 24416 28804 24472 28860
rect 24472 28804 24476 28860
rect 24412 28800 24476 28804
rect 24492 28860 24556 28864
rect 24492 28804 24496 28860
rect 24496 28804 24552 28860
rect 24552 28804 24556 28860
rect 24492 28800 24556 28804
rect 27252 28860 27316 28864
rect 27252 28804 27256 28860
rect 27256 28804 27312 28860
rect 27312 28804 27316 28860
rect 27252 28800 27316 28804
rect 27332 28860 27396 28864
rect 27332 28804 27336 28860
rect 27336 28804 27392 28860
rect 27392 28804 27396 28860
rect 27332 28800 27396 28804
rect 27412 28860 27476 28864
rect 27412 28804 27416 28860
rect 27416 28804 27472 28860
rect 27472 28804 27476 28860
rect 27412 28800 27476 28804
rect 27492 28860 27556 28864
rect 27492 28804 27496 28860
rect 27496 28804 27552 28860
rect 27552 28804 27556 28860
rect 27492 28800 27556 28804
rect 1752 28316 1816 28320
rect 1752 28260 1756 28316
rect 1756 28260 1812 28316
rect 1812 28260 1816 28316
rect 1752 28256 1816 28260
rect 1832 28316 1896 28320
rect 1832 28260 1836 28316
rect 1836 28260 1892 28316
rect 1892 28260 1896 28316
rect 1832 28256 1896 28260
rect 1912 28316 1976 28320
rect 1912 28260 1916 28316
rect 1916 28260 1972 28316
rect 1972 28260 1976 28316
rect 1912 28256 1976 28260
rect 1992 28316 2056 28320
rect 1992 28260 1996 28316
rect 1996 28260 2052 28316
rect 2052 28260 2056 28316
rect 1992 28256 2056 28260
rect 4752 28316 4816 28320
rect 4752 28260 4756 28316
rect 4756 28260 4812 28316
rect 4812 28260 4816 28316
rect 4752 28256 4816 28260
rect 4832 28316 4896 28320
rect 4832 28260 4836 28316
rect 4836 28260 4892 28316
rect 4892 28260 4896 28316
rect 4832 28256 4896 28260
rect 4912 28316 4976 28320
rect 4912 28260 4916 28316
rect 4916 28260 4972 28316
rect 4972 28260 4976 28316
rect 4912 28256 4976 28260
rect 4992 28316 5056 28320
rect 4992 28260 4996 28316
rect 4996 28260 5052 28316
rect 5052 28260 5056 28316
rect 4992 28256 5056 28260
rect 7752 28316 7816 28320
rect 7752 28260 7756 28316
rect 7756 28260 7812 28316
rect 7812 28260 7816 28316
rect 7752 28256 7816 28260
rect 7832 28316 7896 28320
rect 7832 28260 7836 28316
rect 7836 28260 7892 28316
rect 7892 28260 7896 28316
rect 7832 28256 7896 28260
rect 7912 28316 7976 28320
rect 7912 28260 7916 28316
rect 7916 28260 7972 28316
rect 7972 28260 7976 28316
rect 7912 28256 7976 28260
rect 7992 28316 8056 28320
rect 7992 28260 7996 28316
rect 7996 28260 8052 28316
rect 8052 28260 8056 28316
rect 7992 28256 8056 28260
rect 10752 28316 10816 28320
rect 10752 28260 10756 28316
rect 10756 28260 10812 28316
rect 10812 28260 10816 28316
rect 10752 28256 10816 28260
rect 10832 28316 10896 28320
rect 10832 28260 10836 28316
rect 10836 28260 10892 28316
rect 10892 28260 10896 28316
rect 10832 28256 10896 28260
rect 10912 28316 10976 28320
rect 10912 28260 10916 28316
rect 10916 28260 10972 28316
rect 10972 28260 10976 28316
rect 10912 28256 10976 28260
rect 10992 28316 11056 28320
rect 10992 28260 10996 28316
rect 10996 28260 11052 28316
rect 11052 28260 11056 28316
rect 10992 28256 11056 28260
rect 13752 28316 13816 28320
rect 13752 28260 13756 28316
rect 13756 28260 13812 28316
rect 13812 28260 13816 28316
rect 13752 28256 13816 28260
rect 13832 28316 13896 28320
rect 13832 28260 13836 28316
rect 13836 28260 13892 28316
rect 13892 28260 13896 28316
rect 13832 28256 13896 28260
rect 13912 28316 13976 28320
rect 13912 28260 13916 28316
rect 13916 28260 13972 28316
rect 13972 28260 13976 28316
rect 13912 28256 13976 28260
rect 13992 28316 14056 28320
rect 13992 28260 13996 28316
rect 13996 28260 14052 28316
rect 14052 28260 14056 28316
rect 13992 28256 14056 28260
rect 16752 28316 16816 28320
rect 16752 28260 16756 28316
rect 16756 28260 16812 28316
rect 16812 28260 16816 28316
rect 16752 28256 16816 28260
rect 16832 28316 16896 28320
rect 16832 28260 16836 28316
rect 16836 28260 16892 28316
rect 16892 28260 16896 28316
rect 16832 28256 16896 28260
rect 16912 28316 16976 28320
rect 16912 28260 16916 28316
rect 16916 28260 16972 28316
rect 16972 28260 16976 28316
rect 16912 28256 16976 28260
rect 16992 28316 17056 28320
rect 16992 28260 16996 28316
rect 16996 28260 17052 28316
rect 17052 28260 17056 28316
rect 16992 28256 17056 28260
rect 19752 28316 19816 28320
rect 19752 28260 19756 28316
rect 19756 28260 19812 28316
rect 19812 28260 19816 28316
rect 19752 28256 19816 28260
rect 19832 28316 19896 28320
rect 19832 28260 19836 28316
rect 19836 28260 19892 28316
rect 19892 28260 19896 28316
rect 19832 28256 19896 28260
rect 19912 28316 19976 28320
rect 19912 28260 19916 28316
rect 19916 28260 19972 28316
rect 19972 28260 19976 28316
rect 19912 28256 19976 28260
rect 19992 28316 20056 28320
rect 19992 28260 19996 28316
rect 19996 28260 20052 28316
rect 20052 28260 20056 28316
rect 19992 28256 20056 28260
rect 22752 28316 22816 28320
rect 22752 28260 22756 28316
rect 22756 28260 22812 28316
rect 22812 28260 22816 28316
rect 22752 28256 22816 28260
rect 22832 28316 22896 28320
rect 22832 28260 22836 28316
rect 22836 28260 22892 28316
rect 22892 28260 22896 28316
rect 22832 28256 22896 28260
rect 22912 28316 22976 28320
rect 22912 28260 22916 28316
rect 22916 28260 22972 28316
rect 22972 28260 22976 28316
rect 22912 28256 22976 28260
rect 22992 28316 23056 28320
rect 22992 28260 22996 28316
rect 22996 28260 23052 28316
rect 23052 28260 23056 28316
rect 22992 28256 23056 28260
rect 25752 28316 25816 28320
rect 25752 28260 25756 28316
rect 25756 28260 25812 28316
rect 25812 28260 25816 28316
rect 25752 28256 25816 28260
rect 25832 28316 25896 28320
rect 25832 28260 25836 28316
rect 25836 28260 25892 28316
rect 25892 28260 25896 28316
rect 25832 28256 25896 28260
rect 25912 28316 25976 28320
rect 25912 28260 25916 28316
rect 25916 28260 25972 28316
rect 25972 28260 25976 28316
rect 25912 28256 25976 28260
rect 25992 28316 26056 28320
rect 25992 28260 25996 28316
rect 25996 28260 26052 28316
rect 26052 28260 26056 28316
rect 25992 28256 26056 28260
rect 3252 27772 3316 27776
rect 3252 27716 3256 27772
rect 3256 27716 3312 27772
rect 3312 27716 3316 27772
rect 3252 27712 3316 27716
rect 3332 27772 3396 27776
rect 3332 27716 3336 27772
rect 3336 27716 3392 27772
rect 3392 27716 3396 27772
rect 3332 27712 3396 27716
rect 3412 27772 3476 27776
rect 3412 27716 3416 27772
rect 3416 27716 3472 27772
rect 3472 27716 3476 27772
rect 3412 27712 3476 27716
rect 3492 27772 3556 27776
rect 3492 27716 3496 27772
rect 3496 27716 3552 27772
rect 3552 27716 3556 27772
rect 3492 27712 3556 27716
rect 6252 27772 6316 27776
rect 6252 27716 6256 27772
rect 6256 27716 6312 27772
rect 6312 27716 6316 27772
rect 6252 27712 6316 27716
rect 6332 27772 6396 27776
rect 6332 27716 6336 27772
rect 6336 27716 6392 27772
rect 6392 27716 6396 27772
rect 6332 27712 6396 27716
rect 6412 27772 6476 27776
rect 6412 27716 6416 27772
rect 6416 27716 6472 27772
rect 6472 27716 6476 27772
rect 6412 27712 6476 27716
rect 6492 27772 6556 27776
rect 6492 27716 6496 27772
rect 6496 27716 6552 27772
rect 6552 27716 6556 27772
rect 6492 27712 6556 27716
rect 9252 27772 9316 27776
rect 9252 27716 9256 27772
rect 9256 27716 9312 27772
rect 9312 27716 9316 27772
rect 9252 27712 9316 27716
rect 9332 27772 9396 27776
rect 9332 27716 9336 27772
rect 9336 27716 9392 27772
rect 9392 27716 9396 27772
rect 9332 27712 9396 27716
rect 9412 27772 9476 27776
rect 9412 27716 9416 27772
rect 9416 27716 9472 27772
rect 9472 27716 9476 27772
rect 9412 27712 9476 27716
rect 9492 27772 9556 27776
rect 9492 27716 9496 27772
rect 9496 27716 9552 27772
rect 9552 27716 9556 27772
rect 9492 27712 9556 27716
rect 12252 27772 12316 27776
rect 12252 27716 12256 27772
rect 12256 27716 12312 27772
rect 12312 27716 12316 27772
rect 12252 27712 12316 27716
rect 12332 27772 12396 27776
rect 12332 27716 12336 27772
rect 12336 27716 12392 27772
rect 12392 27716 12396 27772
rect 12332 27712 12396 27716
rect 12412 27772 12476 27776
rect 12412 27716 12416 27772
rect 12416 27716 12472 27772
rect 12472 27716 12476 27772
rect 12412 27712 12476 27716
rect 12492 27772 12556 27776
rect 12492 27716 12496 27772
rect 12496 27716 12552 27772
rect 12552 27716 12556 27772
rect 12492 27712 12556 27716
rect 15252 27772 15316 27776
rect 15252 27716 15256 27772
rect 15256 27716 15312 27772
rect 15312 27716 15316 27772
rect 15252 27712 15316 27716
rect 15332 27772 15396 27776
rect 15332 27716 15336 27772
rect 15336 27716 15392 27772
rect 15392 27716 15396 27772
rect 15332 27712 15396 27716
rect 15412 27772 15476 27776
rect 15412 27716 15416 27772
rect 15416 27716 15472 27772
rect 15472 27716 15476 27772
rect 15412 27712 15476 27716
rect 15492 27772 15556 27776
rect 15492 27716 15496 27772
rect 15496 27716 15552 27772
rect 15552 27716 15556 27772
rect 15492 27712 15556 27716
rect 18252 27772 18316 27776
rect 18252 27716 18256 27772
rect 18256 27716 18312 27772
rect 18312 27716 18316 27772
rect 18252 27712 18316 27716
rect 18332 27772 18396 27776
rect 18332 27716 18336 27772
rect 18336 27716 18392 27772
rect 18392 27716 18396 27772
rect 18332 27712 18396 27716
rect 18412 27772 18476 27776
rect 18412 27716 18416 27772
rect 18416 27716 18472 27772
rect 18472 27716 18476 27772
rect 18412 27712 18476 27716
rect 18492 27772 18556 27776
rect 18492 27716 18496 27772
rect 18496 27716 18552 27772
rect 18552 27716 18556 27772
rect 18492 27712 18556 27716
rect 21252 27772 21316 27776
rect 21252 27716 21256 27772
rect 21256 27716 21312 27772
rect 21312 27716 21316 27772
rect 21252 27712 21316 27716
rect 21332 27772 21396 27776
rect 21332 27716 21336 27772
rect 21336 27716 21392 27772
rect 21392 27716 21396 27772
rect 21332 27712 21396 27716
rect 21412 27772 21476 27776
rect 21412 27716 21416 27772
rect 21416 27716 21472 27772
rect 21472 27716 21476 27772
rect 21412 27712 21476 27716
rect 21492 27772 21556 27776
rect 21492 27716 21496 27772
rect 21496 27716 21552 27772
rect 21552 27716 21556 27772
rect 21492 27712 21556 27716
rect 24252 27772 24316 27776
rect 24252 27716 24256 27772
rect 24256 27716 24312 27772
rect 24312 27716 24316 27772
rect 24252 27712 24316 27716
rect 24332 27772 24396 27776
rect 24332 27716 24336 27772
rect 24336 27716 24392 27772
rect 24392 27716 24396 27772
rect 24332 27712 24396 27716
rect 24412 27772 24476 27776
rect 24412 27716 24416 27772
rect 24416 27716 24472 27772
rect 24472 27716 24476 27772
rect 24412 27712 24476 27716
rect 24492 27772 24556 27776
rect 24492 27716 24496 27772
rect 24496 27716 24552 27772
rect 24552 27716 24556 27772
rect 24492 27712 24556 27716
rect 27252 27772 27316 27776
rect 27252 27716 27256 27772
rect 27256 27716 27312 27772
rect 27312 27716 27316 27772
rect 27252 27712 27316 27716
rect 27332 27772 27396 27776
rect 27332 27716 27336 27772
rect 27336 27716 27392 27772
rect 27392 27716 27396 27772
rect 27332 27712 27396 27716
rect 27412 27772 27476 27776
rect 27412 27716 27416 27772
rect 27416 27716 27472 27772
rect 27472 27716 27476 27772
rect 27412 27712 27476 27716
rect 27492 27772 27556 27776
rect 27492 27716 27496 27772
rect 27496 27716 27552 27772
rect 27552 27716 27556 27772
rect 27492 27712 27556 27716
rect 1752 27228 1816 27232
rect 1752 27172 1756 27228
rect 1756 27172 1812 27228
rect 1812 27172 1816 27228
rect 1752 27168 1816 27172
rect 1832 27228 1896 27232
rect 1832 27172 1836 27228
rect 1836 27172 1892 27228
rect 1892 27172 1896 27228
rect 1832 27168 1896 27172
rect 1912 27228 1976 27232
rect 1912 27172 1916 27228
rect 1916 27172 1972 27228
rect 1972 27172 1976 27228
rect 1912 27168 1976 27172
rect 1992 27228 2056 27232
rect 1992 27172 1996 27228
rect 1996 27172 2052 27228
rect 2052 27172 2056 27228
rect 1992 27168 2056 27172
rect 4752 27228 4816 27232
rect 4752 27172 4756 27228
rect 4756 27172 4812 27228
rect 4812 27172 4816 27228
rect 4752 27168 4816 27172
rect 4832 27228 4896 27232
rect 4832 27172 4836 27228
rect 4836 27172 4892 27228
rect 4892 27172 4896 27228
rect 4832 27168 4896 27172
rect 4912 27228 4976 27232
rect 4912 27172 4916 27228
rect 4916 27172 4972 27228
rect 4972 27172 4976 27228
rect 4912 27168 4976 27172
rect 4992 27228 5056 27232
rect 4992 27172 4996 27228
rect 4996 27172 5052 27228
rect 5052 27172 5056 27228
rect 4992 27168 5056 27172
rect 7752 27228 7816 27232
rect 7752 27172 7756 27228
rect 7756 27172 7812 27228
rect 7812 27172 7816 27228
rect 7752 27168 7816 27172
rect 7832 27228 7896 27232
rect 7832 27172 7836 27228
rect 7836 27172 7892 27228
rect 7892 27172 7896 27228
rect 7832 27168 7896 27172
rect 7912 27228 7976 27232
rect 7912 27172 7916 27228
rect 7916 27172 7972 27228
rect 7972 27172 7976 27228
rect 7912 27168 7976 27172
rect 7992 27228 8056 27232
rect 7992 27172 7996 27228
rect 7996 27172 8052 27228
rect 8052 27172 8056 27228
rect 7992 27168 8056 27172
rect 10752 27228 10816 27232
rect 10752 27172 10756 27228
rect 10756 27172 10812 27228
rect 10812 27172 10816 27228
rect 10752 27168 10816 27172
rect 10832 27228 10896 27232
rect 10832 27172 10836 27228
rect 10836 27172 10892 27228
rect 10892 27172 10896 27228
rect 10832 27168 10896 27172
rect 10912 27228 10976 27232
rect 10912 27172 10916 27228
rect 10916 27172 10972 27228
rect 10972 27172 10976 27228
rect 10912 27168 10976 27172
rect 10992 27228 11056 27232
rect 10992 27172 10996 27228
rect 10996 27172 11052 27228
rect 11052 27172 11056 27228
rect 10992 27168 11056 27172
rect 13752 27228 13816 27232
rect 13752 27172 13756 27228
rect 13756 27172 13812 27228
rect 13812 27172 13816 27228
rect 13752 27168 13816 27172
rect 13832 27228 13896 27232
rect 13832 27172 13836 27228
rect 13836 27172 13892 27228
rect 13892 27172 13896 27228
rect 13832 27168 13896 27172
rect 13912 27228 13976 27232
rect 13912 27172 13916 27228
rect 13916 27172 13972 27228
rect 13972 27172 13976 27228
rect 13912 27168 13976 27172
rect 13992 27228 14056 27232
rect 13992 27172 13996 27228
rect 13996 27172 14052 27228
rect 14052 27172 14056 27228
rect 13992 27168 14056 27172
rect 16752 27228 16816 27232
rect 16752 27172 16756 27228
rect 16756 27172 16812 27228
rect 16812 27172 16816 27228
rect 16752 27168 16816 27172
rect 16832 27228 16896 27232
rect 16832 27172 16836 27228
rect 16836 27172 16892 27228
rect 16892 27172 16896 27228
rect 16832 27168 16896 27172
rect 16912 27228 16976 27232
rect 16912 27172 16916 27228
rect 16916 27172 16972 27228
rect 16972 27172 16976 27228
rect 16912 27168 16976 27172
rect 16992 27228 17056 27232
rect 16992 27172 16996 27228
rect 16996 27172 17052 27228
rect 17052 27172 17056 27228
rect 16992 27168 17056 27172
rect 19752 27228 19816 27232
rect 19752 27172 19756 27228
rect 19756 27172 19812 27228
rect 19812 27172 19816 27228
rect 19752 27168 19816 27172
rect 19832 27228 19896 27232
rect 19832 27172 19836 27228
rect 19836 27172 19892 27228
rect 19892 27172 19896 27228
rect 19832 27168 19896 27172
rect 19912 27228 19976 27232
rect 19912 27172 19916 27228
rect 19916 27172 19972 27228
rect 19972 27172 19976 27228
rect 19912 27168 19976 27172
rect 19992 27228 20056 27232
rect 19992 27172 19996 27228
rect 19996 27172 20052 27228
rect 20052 27172 20056 27228
rect 19992 27168 20056 27172
rect 22752 27228 22816 27232
rect 22752 27172 22756 27228
rect 22756 27172 22812 27228
rect 22812 27172 22816 27228
rect 22752 27168 22816 27172
rect 22832 27228 22896 27232
rect 22832 27172 22836 27228
rect 22836 27172 22892 27228
rect 22892 27172 22896 27228
rect 22832 27168 22896 27172
rect 22912 27228 22976 27232
rect 22912 27172 22916 27228
rect 22916 27172 22972 27228
rect 22972 27172 22976 27228
rect 22912 27168 22976 27172
rect 22992 27228 23056 27232
rect 22992 27172 22996 27228
rect 22996 27172 23052 27228
rect 23052 27172 23056 27228
rect 22992 27168 23056 27172
rect 25752 27228 25816 27232
rect 25752 27172 25756 27228
rect 25756 27172 25812 27228
rect 25812 27172 25816 27228
rect 25752 27168 25816 27172
rect 25832 27228 25896 27232
rect 25832 27172 25836 27228
rect 25836 27172 25892 27228
rect 25892 27172 25896 27228
rect 25832 27168 25896 27172
rect 25912 27228 25976 27232
rect 25912 27172 25916 27228
rect 25916 27172 25972 27228
rect 25972 27172 25976 27228
rect 25912 27168 25976 27172
rect 25992 27228 26056 27232
rect 25992 27172 25996 27228
rect 25996 27172 26052 27228
rect 26052 27172 26056 27228
rect 25992 27168 26056 27172
rect 3252 26684 3316 26688
rect 3252 26628 3256 26684
rect 3256 26628 3312 26684
rect 3312 26628 3316 26684
rect 3252 26624 3316 26628
rect 3332 26684 3396 26688
rect 3332 26628 3336 26684
rect 3336 26628 3392 26684
rect 3392 26628 3396 26684
rect 3332 26624 3396 26628
rect 3412 26684 3476 26688
rect 3412 26628 3416 26684
rect 3416 26628 3472 26684
rect 3472 26628 3476 26684
rect 3412 26624 3476 26628
rect 3492 26684 3556 26688
rect 3492 26628 3496 26684
rect 3496 26628 3552 26684
rect 3552 26628 3556 26684
rect 3492 26624 3556 26628
rect 6252 26684 6316 26688
rect 6252 26628 6256 26684
rect 6256 26628 6312 26684
rect 6312 26628 6316 26684
rect 6252 26624 6316 26628
rect 6332 26684 6396 26688
rect 6332 26628 6336 26684
rect 6336 26628 6392 26684
rect 6392 26628 6396 26684
rect 6332 26624 6396 26628
rect 6412 26684 6476 26688
rect 6412 26628 6416 26684
rect 6416 26628 6472 26684
rect 6472 26628 6476 26684
rect 6412 26624 6476 26628
rect 6492 26684 6556 26688
rect 6492 26628 6496 26684
rect 6496 26628 6552 26684
rect 6552 26628 6556 26684
rect 6492 26624 6556 26628
rect 9252 26684 9316 26688
rect 9252 26628 9256 26684
rect 9256 26628 9312 26684
rect 9312 26628 9316 26684
rect 9252 26624 9316 26628
rect 9332 26684 9396 26688
rect 9332 26628 9336 26684
rect 9336 26628 9392 26684
rect 9392 26628 9396 26684
rect 9332 26624 9396 26628
rect 9412 26684 9476 26688
rect 9412 26628 9416 26684
rect 9416 26628 9472 26684
rect 9472 26628 9476 26684
rect 9412 26624 9476 26628
rect 9492 26684 9556 26688
rect 9492 26628 9496 26684
rect 9496 26628 9552 26684
rect 9552 26628 9556 26684
rect 9492 26624 9556 26628
rect 12252 26684 12316 26688
rect 12252 26628 12256 26684
rect 12256 26628 12312 26684
rect 12312 26628 12316 26684
rect 12252 26624 12316 26628
rect 12332 26684 12396 26688
rect 12332 26628 12336 26684
rect 12336 26628 12392 26684
rect 12392 26628 12396 26684
rect 12332 26624 12396 26628
rect 12412 26684 12476 26688
rect 12412 26628 12416 26684
rect 12416 26628 12472 26684
rect 12472 26628 12476 26684
rect 12412 26624 12476 26628
rect 12492 26684 12556 26688
rect 12492 26628 12496 26684
rect 12496 26628 12552 26684
rect 12552 26628 12556 26684
rect 12492 26624 12556 26628
rect 15252 26684 15316 26688
rect 15252 26628 15256 26684
rect 15256 26628 15312 26684
rect 15312 26628 15316 26684
rect 15252 26624 15316 26628
rect 15332 26684 15396 26688
rect 15332 26628 15336 26684
rect 15336 26628 15392 26684
rect 15392 26628 15396 26684
rect 15332 26624 15396 26628
rect 15412 26684 15476 26688
rect 15412 26628 15416 26684
rect 15416 26628 15472 26684
rect 15472 26628 15476 26684
rect 15412 26624 15476 26628
rect 15492 26684 15556 26688
rect 15492 26628 15496 26684
rect 15496 26628 15552 26684
rect 15552 26628 15556 26684
rect 15492 26624 15556 26628
rect 18252 26684 18316 26688
rect 18252 26628 18256 26684
rect 18256 26628 18312 26684
rect 18312 26628 18316 26684
rect 18252 26624 18316 26628
rect 18332 26684 18396 26688
rect 18332 26628 18336 26684
rect 18336 26628 18392 26684
rect 18392 26628 18396 26684
rect 18332 26624 18396 26628
rect 18412 26684 18476 26688
rect 18412 26628 18416 26684
rect 18416 26628 18472 26684
rect 18472 26628 18476 26684
rect 18412 26624 18476 26628
rect 18492 26684 18556 26688
rect 18492 26628 18496 26684
rect 18496 26628 18552 26684
rect 18552 26628 18556 26684
rect 18492 26624 18556 26628
rect 21252 26684 21316 26688
rect 21252 26628 21256 26684
rect 21256 26628 21312 26684
rect 21312 26628 21316 26684
rect 21252 26624 21316 26628
rect 21332 26684 21396 26688
rect 21332 26628 21336 26684
rect 21336 26628 21392 26684
rect 21392 26628 21396 26684
rect 21332 26624 21396 26628
rect 21412 26684 21476 26688
rect 21412 26628 21416 26684
rect 21416 26628 21472 26684
rect 21472 26628 21476 26684
rect 21412 26624 21476 26628
rect 21492 26684 21556 26688
rect 21492 26628 21496 26684
rect 21496 26628 21552 26684
rect 21552 26628 21556 26684
rect 21492 26624 21556 26628
rect 24252 26684 24316 26688
rect 24252 26628 24256 26684
rect 24256 26628 24312 26684
rect 24312 26628 24316 26684
rect 24252 26624 24316 26628
rect 24332 26684 24396 26688
rect 24332 26628 24336 26684
rect 24336 26628 24392 26684
rect 24392 26628 24396 26684
rect 24332 26624 24396 26628
rect 24412 26684 24476 26688
rect 24412 26628 24416 26684
rect 24416 26628 24472 26684
rect 24472 26628 24476 26684
rect 24412 26624 24476 26628
rect 24492 26684 24556 26688
rect 24492 26628 24496 26684
rect 24496 26628 24552 26684
rect 24552 26628 24556 26684
rect 24492 26624 24556 26628
rect 27252 26684 27316 26688
rect 27252 26628 27256 26684
rect 27256 26628 27312 26684
rect 27312 26628 27316 26684
rect 27252 26624 27316 26628
rect 27332 26684 27396 26688
rect 27332 26628 27336 26684
rect 27336 26628 27392 26684
rect 27392 26628 27396 26684
rect 27332 26624 27396 26628
rect 27412 26684 27476 26688
rect 27412 26628 27416 26684
rect 27416 26628 27472 26684
rect 27472 26628 27476 26684
rect 27412 26624 27476 26628
rect 27492 26684 27556 26688
rect 27492 26628 27496 26684
rect 27496 26628 27552 26684
rect 27552 26628 27556 26684
rect 27492 26624 27556 26628
rect 1752 26140 1816 26144
rect 1752 26084 1756 26140
rect 1756 26084 1812 26140
rect 1812 26084 1816 26140
rect 1752 26080 1816 26084
rect 1832 26140 1896 26144
rect 1832 26084 1836 26140
rect 1836 26084 1892 26140
rect 1892 26084 1896 26140
rect 1832 26080 1896 26084
rect 1912 26140 1976 26144
rect 1912 26084 1916 26140
rect 1916 26084 1972 26140
rect 1972 26084 1976 26140
rect 1912 26080 1976 26084
rect 1992 26140 2056 26144
rect 1992 26084 1996 26140
rect 1996 26084 2052 26140
rect 2052 26084 2056 26140
rect 1992 26080 2056 26084
rect 4752 26140 4816 26144
rect 4752 26084 4756 26140
rect 4756 26084 4812 26140
rect 4812 26084 4816 26140
rect 4752 26080 4816 26084
rect 4832 26140 4896 26144
rect 4832 26084 4836 26140
rect 4836 26084 4892 26140
rect 4892 26084 4896 26140
rect 4832 26080 4896 26084
rect 4912 26140 4976 26144
rect 4912 26084 4916 26140
rect 4916 26084 4972 26140
rect 4972 26084 4976 26140
rect 4912 26080 4976 26084
rect 4992 26140 5056 26144
rect 4992 26084 4996 26140
rect 4996 26084 5052 26140
rect 5052 26084 5056 26140
rect 4992 26080 5056 26084
rect 7752 26140 7816 26144
rect 7752 26084 7756 26140
rect 7756 26084 7812 26140
rect 7812 26084 7816 26140
rect 7752 26080 7816 26084
rect 7832 26140 7896 26144
rect 7832 26084 7836 26140
rect 7836 26084 7892 26140
rect 7892 26084 7896 26140
rect 7832 26080 7896 26084
rect 7912 26140 7976 26144
rect 7912 26084 7916 26140
rect 7916 26084 7972 26140
rect 7972 26084 7976 26140
rect 7912 26080 7976 26084
rect 7992 26140 8056 26144
rect 7992 26084 7996 26140
rect 7996 26084 8052 26140
rect 8052 26084 8056 26140
rect 7992 26080 8056 26084
rect 10752 26140 10816 26144
rect 10752 26084 10756 26140
rect 10756 26084 10812 26140
rect 10812 26084 10816 26140
rect 10752 26080 10816 26084
rect 10832 26140 10896 26144
rect 10832 26084 10836 26140
rect 10836 26084 10892 26140
rect 10892 26084 10896 26140
rect 10832 26080 10896 26084
rect 10912 26140 10976 26144
rect 10912 26084 10916 26140
rect 10916 26084 10972 26140
rect 10972 26084 10976 26140
rect 10912 26080 10976 26084
rect 10992 26140 11056 26144
rect 10992 26084 10996 26140
rect 10996 26084 11052 26140
rect 11052 26084 11056 26140
rect 10992 26080 11056 26084
rect 13752 26140 13816 26144
rect 13752 26084 13756 26140
rect 13756 26084 13812 26140
rect 13812 26084 13816 26140
rect 13752 26080 13816 26084
rect 13832 26140 13896 26144
rect 13832 26084 13836 26140
rect 13836 26084 13892 26140
rect 13892 26084 13896 26140
rect 13832 26080 13896 26084
rect 13912 26140 13976 26144
rect 13912 26084 13916 26140
rect 13916 26084 13972 26140
rect 13972 26084 13976 26140
rect 13912 26080 13976 26084
rect 13992 26140 14056 26144
rect 13992 26084 13996 26140
rect 13996 26084 14052 26140
rect 14052 26084 14056 26140
rect 13992 26080 14056 26084
rect 16752 26140 16816 26144
rect 16752 26084 16756 26140
rect 16756 26084 16812 26140
rect 16812 26084 16816 26140
rect 16752 26080 16816 26084
rect 16832 26140 16896 26144
rect 16832 26084 16836 26140
rect 16836 26084 16892 26140
rect 16892 26084 16896 26140
rect 16832 26080 16896 26084
rect 16912 26140 16976 26144
rect 16912 26084 16916 26140
rect 16916 26084 16972 26140
rect 16972 26084 16976 26140
rect 16912 26080 16976 26084
rect 16992 26140 17056 26144
rect 16992 26084 16996 26140
rect 16996 26084 17052 26140
rect 17052 26084 17056 26140
rect 16992 26080 17056 26084
rect 19752 26140 19816 26144
rect 19752 26084 19756 26140
rect 19756 26084 19812 26140
rect 19812 26084 19816 26140
rect 19752 26080 19816 26084
rect 19832 26140 19896 26144
rect 19832 26084 19836 26140
rect 19836 26084 19892 26140
rect 19892 26084 19896 26140
rect 19832 26080 19896 26084
rect 19912 26140 19976 26144
rect 19912 26084 19916 26140
rect 19916 26084 19972 26140
rect 19972 26084 19976 26140
rect 19912 26080 19976 26084
rect 19992 26140 20056 26144
rect 19992 26084 19996 26140
rect 19996 26084 20052 26140
rect 20052 26084 20056 26140
rect 19992 26080 20056 26084
rect 22752 26140 22816 26144
rect 22752 26084 22756 26140
rect 22756 26084 22812 26140
rect 22812 26084 22816 26140
rect 22752 26080 22816 26084
rect 22832 26140 22896 26144
rect 22832 26084 22836 26140
rect 22836 26084 22892 26140
rect 22892 26084 22896 26140
rect 22832 26080 22896 26084
rect 22912 26140 22976 26144
rect 22912 26084 22916 26140
rect 22916 26084 22972 26140
rect 22972 26084 22976 26140
rect 22912 26080 22976 26084
rect 22992 26140 23056 26144
rect 22992 26084 22996 26140
rect 22996 26084 23052 26140
rect 23052 26084 23056 26140
rect 22992 26080 23056 26084
rect 25752 26140 25816 26144
rect 25752 26084 25756 26140
rect 25756 26084 25812 26140
rect 25812 26084 25816 26140
rect 25752 26080 25816 26084
rect 25832 26140 25896 26144
rect 25832 26084 25836 26140
rect 25836 26084 25892 26140
rect 25892 26084 25896 26140
rect 25832 26080 25896 26084
rect 25912 26140 25976 26144
rect 25912 26084 25916 26140
rect 25916 26084 25972 26140
rect 25972 26084 25976 26140
rect 25912 26080 25976 26084
rect 25992 26140 26056 26144
rect 25992 26084 25996 26140
rect 25996 26084 26052 26140
rect 26052 26084 26056 26140
rect 25992 26080 26056 26084
rect 3252 25596 3316 25600
rect 3252 25540 3256 25596
rect 3256 25540 3312 25596
rect 3312 25540 3316 25596
rect 3252 25536 3316 25540
rect 3332 25596 3396 25600
rect 3332 25540 3336 25596
rect 3336 25540 3392 25596
rect 3392 25540 3396 25596
rect 3332 25536 3396 25540
rect 3412 25596 3476 25600
rect 3412 25540 3416 25596
rect 3416 25540 3472 25596
rect 3472 25540 3476 25596
rect 3412 25536 3476 25540
rect 3492 25596 3556 25600
rect 3492 25540 3496 25596
rect 3496 25540 3552 25596
rect 3552 25540 3556 25596
rect 3492 25536 3556 25540
rect 6252 25596 6316 25600
rect 6252 25540 6256 25596
rect 6256 25540 6312 25596
rect 6312 25540 6316 25596
rect 6252 25536 6316 25540
rect 6332 25596 6396 25600
rect 6332 25540 6336 25596
rect 6336 25540 6392 25596
rect 6392 25540 6396 25596
rect 6332 25536 6396 25540
rect 6412 25596 6476 25600
rect 6412 25540 6416 25596
rect 6416 25540 6472 25596
rect 6472 25540 6476 25596
rect 6412 25536 6476 25540
rect 6492 25596 6556 25600
rect 6492 25540 6496 25596
rect 6496 25540 6552 25596
rect 6552 25540 6556 25596
rect 6492 25536 6556 25540
rect 9252 25596 9316 25600
rect 9252 25540 9256 25596
rect 9256 25540 9312 25596
rect 9312 25540 9316 25596
rect 9252 25536 9316 25540
rect 9332 25596 9396 25600
rect 9332 25540 9336 25596
rect 9336 25540 9392 25596
rect 9392 25540 9396 25596
rect 9332 25536 9396 25540
rect 9412 25596 9476 25600
rect 9412 25540 9416 25596
rect 9416 25540 9472 25596
rect 9472 25540 9476 25596
rect 9412 25536 9476 25540
rect 9492 25596 9556 25600
rect 9492 25540 9496 25596
rect 9496 25540 9552 25596
rect 9552 25540 9556 25596
rect 9492 25536 9556 25540
rect 12252 25596 12316 25600
rect 12252 25540 12256 25596
rect 12256 25540 12312 25596
rect 12312 25540 12316 25596
rect 12252 25536 12316 25540
rect 12332 25596 12396 25600
rect 12332 25540 12336 25596
rect 12336 25540 12392 25596
rect 12392 25540 12396 25596
rect 12332 25536 12396 25540
rect 12412 25596 12476 25600
rect 12412 25540 12416 25596
rect 12416 25540 12472 25596
rect 12472 25540 12476 25596
rect 12412 25536 12476 25540
rect 12492 25596 12556 25600
rect 12492 25540 12496 25596
rect 12496 25540 12552 25596
rect 12552 25540 12556 25596
rect 12492 25536 12556 25540
rect 15252 25596 15316 25600
rect 15252 25540 15256 25596
rect 15256 25540 15312 25596
rect 15312 25540 15316 25596
rect 15252 25536 15316 25540
rect 15332 25596 15396 25600
rect 15332 25540 15336 25596
rect 15336 25540 15392 25596
rect 15392 25540 15396 25596
rect 15332 25536 15396 25540
rect 15412 25596 15476 25600
rect 15412 25540 15416 25596
rect 15416 25540 15472 25596
rect 15472 25540 15476 25596
rect 15412 25536 15476 25540
rect 15492 25596 15556 25600
rect 15492 25540 15496 25596
rect 15496 25540 15552 25596
rect 15552 25540 15556 25596
rect 15492 25536 15556 25540
rect 18252 25596 18316 25600
rect 18252 25540 18256 25596
rect 18256 25540 18312 25596
rect 18312 25540 18316 25596
rect 18252 25536 18316 25540
rect 18332 25596 18396 25600
rect 18332 25540 18336 25596
rect 18336 25540 18392 25596
rect 18392 25540 18396 25596
rect 18332 25536 18396 25540
rect 18412 25596 18476 25600
rect 18412 25540 18416 25596
rect 18416 25540 18472 25596
rect 18472 25540 18476 25596
rect 18412 25536 18476 25540
rect 18492 25596 18556 25600
rect 18492 25540 18496 25596
rect 18496 25540 18552 25596
rect 18552 25540 18556 25596
rect 18492 25536 18556 25540
rect 21252 25596 21316 25600
rect 21252 25540 21256 25596
rect 21256 25540 21312 25596
rect 21312 25540 21316 25596
rect 21252 25536 21316 25540
rect 21332 25596 21396 25600
rect 21332 25540 21336 25596
rect 21336 25540 21392 25596
rect 21392 25540 21396 25596
rect 21332 25536 21396 25540
rect 21412 25596 21476 25600
rect 21412 25540 21416 25596
rect 21416 25540 21472 25596
rect 21472 25540 21476 25596
rect 21412 25536 21476 25540
rect 21492 25596 21556 25600
rect 21492 25540 21496 25596
rect 21496 25540 21552 25596
rect 21552 25540 21556 25596
rect 21492 25536 21556 25540
rect 24252 25596 24316 25600
rect 24252 25540 24256 25596
rect 24256 25540 24312 25596
rect 24312 25540 24316 25596
rect 24252 25536 24316 25540
rect 24332 25596 24396 25600
rect 24332 25540 24336 25596
rect 24336 25540 24392 25596
rect 24392 25540 24396 25596
rect 24332 25536 24396 25540
rect 24412 25596 24476 25600
rect 24412 25540 24416 25596
rect 24416 25540 24472 25596
rect 24472 25540 24476 25596
rect 24412 25536 24476 25540
rect 24492 25596 24556 25600
rect 24492 25540 24496 25596
rect 24496 25540 24552 25596
rect 24552 25540 24556 25596
rect 24492 25536 24556 25540
rect 27252 25596 27316 25600
rect 27252 25540 27256 25596
rect 27256 25540 27312 25596
rect 27312 25540 27316 25596
rect 27252 25536 27316 25540
rect 27332 25596 27396 25600
rect 27332 25540 27336 25596
rect 27336 25540 27392 25596
rect 27392 25540 27396 25596
rect 27332 25536 27396 25540
rect 27412 25596 27476 25600
rect 27412 25540 27416 25596
rect 27416 25540 27472 25596
rect 27472 25540 27476 25596
rect 27412 25536 27476 25540
rect 27492 25596 27556 25600
rect 27492 25540 27496 25596
rect 27496 25540 27552 25596
rect 27552 25540 27556 25596
rect 27492 25536 27556 25540
rect 1752 25052 1816 25056
rect 1752 24996 1756 25052
rect 1756 24996 1812 25052
rect 1812 24996 1816 25052
rect 1752 24992 1816 24996
rect 1832 25052 1896 25056
rect 1832 24996 1836 25052
rect 1836 24996 1892 25052
rect 1892 24996 1896 25052
rect 1832 24992 1896 24996
rect 1912 25052 1976 25056
rect 1912 24996 1916 25052
rect 1916 24996 1972 25052
rect 1972 24996 1976 25052
rect 1912 24992 1976 24996
rect 1992 25052 2056 25056
rect 1992 24996 1996 25052
rect 1996 24996 2052 25052
rect 2052 24996 2056 25052
rect 1992 24992 2056 24996
rect 4752 25052 4816 25056
rect 4752 24996 4756 25052
rect 4756 24996 4812 25052
rect 4812 24996 4816 25052
rect 4752 24992 4816 24996
rect 4832 25052 4896 25056
rect 4832 24996 4836 25052
rect 4836 24996 4892 25052
rect 4892 24996 4896 25052
rect 4832 24992 4896 24996
rect 4912 25052 4976 25056
rect 4912 24996 4916 25052
rect 4916 24996 4972 25052
rect 4972 24996 4976 25052
rect 4912 24992 4976 24996
rect 4992 25052 5056 25056
rect 4992 24996 4996 25052
rect 4996 24996 5052 25052
rect 5052 24996 5056 25052
rect 4992 24992 5056 24996
rect 7752 25052 7816 25056
rect 7752 24996 7756 25052
rect 7756 24996 7812 25052
rect 7812 24996 7816 25052
rect 7752 24992 7816 24996
rect 7832 25052 7896 25056
rect 7832 24996 7836 25052
rect 7836 24996 7892 25052
rect 7892 24996 7896 25052
rect 7832 24992 7896 24996
rect 7912 25052 7976 25056
rect 7912 24996 7916 25052
rect 7916 24996 7972 25052
rect 7972 24996 7976 25052
rect 7912 24992 7976 24996
rect 7992 25052 8056 25056
rect 7992 24996 7996 25052
rect 7996 24996 8052 25052
rect 8052 24996 8056 25052
rect 7992 24992 8056 24996
rect 10752 25052 10816 25056
rect 10752 24996 10756 25052
rect 10756 24996 10812 25052
rect 10812 24996 10816 25052
rect 10752 24992 10816 24996
rect 10832 25052 10896 25056
rect 10832 24996 10836 25052
rect 10836 24996 10892 25052
rect 10892 24996 10896 25052
rect 10832 24992 10896 24996
rect 10912 25052 10976 25056
rect 10912 24996 10916 25052
rect 10916 24996 10972 25052
rect 10972 24996 10976 25052
rect 10912 24992 10976 24996
rect 10992 25052 11056 25056
rect 10992 24996 10996 25052
rect 10996 24996 11052 25052
rect 11052 24996 11056 25052
rect 10992 24992 11056 24996
rect 13752 25052 13816 25056
rect 13752 24996 13756 25052
rect 13756 24996 13812 25052
rect 13812 24996 13816 25052
rect 13752 24992 13816 24996
rect 13832 25052 13896 25056
rect 13832 24996 13836 25052
rect 13836 24996 13892 25052
rect 13892 24996 13896 25052
rect 13832 24992 13896 24996
rect 13912 25052 13976 25056
rect 13912 24996 13916 25052
rect 13916 24996 13972 25052
rect 13972 24996 13976 25052
rect 13912 24992 13976 24996
rect 13992 25052 14056 25056
rect 13992 24996 13996 25052
rect 13996 24996 14052 25052
rect 14052 24996 14056 25052
rect 13992 24992 14056 24996
rect 16752 25052 16816 25056
rect 16752 24996 16756 25052
rect 16756 24996 16812 25052
rect 16812 24996 16816 25052
rect 16752 24992 16816 24996
rect 16832 25052 16896 25056
rect 16832 24996 16836 25052
rect 16836 24996 16892 25052
rect 16892 24996 16896 25052
rect 16832 24992 16896 24996
rect 16912 25052 16976 25056
rect 16912 24996 16916 25052
rect 16916 24996 16972 25052
rect 16972 24996 16976 25052
rect 16912 24992 16976 24996
rect 16992 25052 17056 25056
rect 16992 24996 16996 25052
rect 16996 24996 17052 25052
rect 17052 24996 17056 25052
rect 16992 24992 17056 24996
rect 19752 25052 19816 25056
rect 19752 24996 19756 25052
rect 19756 24996 19812 25052
rect 19812 24996 19816 25052
rect 19752 24992 19816 24996
rect 19832 25052 19896 25056
rect 19832 24996 19836 25052
rect 19836 24996 19892 25052
rect 19892 24996 19896 25052
rect 19832 24992 19896 24996
rect 19912 25052 19976 25056
rect 19912 24996 19916 25052
rect 19916 24996 19972 25052
rect 19972 24996 19976 25052
rect 19912 24992 19976 24996
rect 19992 25052 20056 25056
rect 19992 24996 19996 25052
rect 19996 24996 20052 25052
rect 20052 24996 20056 25052
rect 19992 24992 20056 24996
rect 22752 25052 22816 25056
rect 22752 24996 22756 25052
rect 22756 24996 22812 25052
rect 22812 24996 22816 25052
rect 22752 24992 22816 24996
rect 22832 25052 22896 25056
rect 22832 24996 22836 25052
rect 22836 24996 22892 25052
rect 22892 24996 22896 25052
rect 22832 24992 22896 24996
rect 22912 25052 22976 25056
rect 22912 24996 22916 25052
rect 22916 24996 22972 25052
rect 22972 24996 22976 25052
rect 22912 24992 22976 24996
rect 22992 25052 23056 25056
rect 22992 24996 22996 25052
rect 22996 24996 23052 25052
rect 23052 24996 23056 25052
rect 22992 24992 23056 24996
rect 25752 25052 25816 25056
rect 25752 24996 25756 25052
rect 25756 24996 25812 25052
rect 25812 24996 25816 25052
rect 25752 24992 25816 24996
rect 25832 25052 25896 25056
rect 25832 24996 25836 25052
rect 25836 24996 25892 25052
rect 25892 24996 25896 25052
rect 25832 24992 25896 24996
rect 25912 25052 25976 25056
rect 25912 24996 25916 25052
rect 25916 24996 25972 25052
rect 25972 24996 25976 25052
rect 25912 24992 25976 24996
rect 25992 25052 26056 25056
rect 25992 24996 25996 25052
rect 25996 24996 26052 25052
rect 26052 24996 26056 25052
rect 25992 24992 26056 24996
rect 3252 24508 3316 24512
rect 3252 24452 3256 24508
rect 3256 24452 3312 24508
rect 3312 24452 3316 24508
rect 3252 24448 3316 24452
rect 3332 24508 3396 24512
rect 3332 24452 3336 24508
rect 3336 24452 3392 24508
rect 3392 24452 3396 24508
rect 3332 24448 3396 24452
rect 3412 24508 3476 24512
rect 3412 24452 3416 24508
rect 3416 24452 3472 24508
rect 3472 24452 3476 24508
rect 3412 24448 3476 24452
rect 3492 24508 3556 24512
rect 3492 24452 3496 24508
rect 3496 24452 3552 24508
rect 3552 24452 3556 24508
rect 3492 24448 3556 24452
rect 6252 24508 6316 24512
rect 6252 24452 6256 24508
rect 6256 24452 6312 24508
rect 6312 24452 6316 24508
rect 6252 24448 6316 24452
rect 6332 24508 6396 24512
rect 6332 24452 6336 24508
rect 6336 24452 6392 24508
rect 6392 24452 6396 24508
rect 6332 24448 6396 24452
rect 6412 24508 6476 24512
rect 6412 24452 6416 24508
rect 6416 24452 6472 24508
rect 6472 24452 6476 24508
rect 6412 24448 6476 24452
rect 6492 24508 6556 24512
rect 6492 24452 6496 24508
rect 6496 24452 6552 24508
rect 6552 24452 6556 24508
rect 6492 24448 6556 24452
rect 9252 24508 9316 24512
rect 9252 24452 9256 24508
rect 9256 24452 9312 24508
rect 9312 24452 9316 24508
rect 9252 24448 9316 24452
rect 9332 24508 9396 24512
rect 9332 24452 9336 24508
rect 9336 24452 9392 24508
rect 9392 24452 9396 24508
rect 9332 24448 9396 24452
rect 9412 24508 9476 24512
rect 9412 24452 9416 24508
rect 9416 24452 9472 24508
rect 9472 24452 9476 24508
rect 9412 24448 9476 24452
rect 9492 24508 9556 24512
rect 9492 24452 9496 24508
rect 9496 24452 9552 24508
rect 9552 24452 9556 24508
rect 9492 24448 9556 24452
rect 12252 24508 12316 24512
rect 12252 24452 12256 24508
rect 12256 24452 12312 24508
rect 12312 24452 12316 24508
rect 12252 24448 12316 24452
rect 12332 24508 12396 24512
rect 12332 24452 12336 24508
rect 12336 24452 12392 24508
rect 12392 24452 12396 24508
rect 12332 24448 12396 24452
rect 12412 24508 12476 24512
rect 12412 24452 12416 24508
rect 12416 24452 12472 24508
rect 12472 24452 12476 24508
rect 12412 24448 12476 24452
rect 12492 24508 12556 24512
rect 12492 24452 12496 24508
rect 12496 24452 12552 24508
rect 12552 24452 12556 24508
rect 12492 24448 12556 24452
rect 15252 24508 15316 24512
rect 15252 24452 15256 24508
rect 15256 24452 15312 24508
rect 15312 24452 15316 24508
rect 15252 24448 15316 24452
rect 15332 24508 15396 24512
rect 15332 24452 15336 24508
rect 15336 24452 15392 24508
rect 15392 24452 15396 24508
rect 15332 24448 15396 24452
rect 15412 24508 15476 24512
rect 15412 24452 15416 24508
rect 15416 24452 15472 24508
rect 15472 24452 15476 24508
rect 15412 24448 15476 24452
rect 15492 24508 15556 24512
rect 15492 24452 15496 24508
rect 15496 24452 15552 24508
rect 15552 24452 15556 24508
rect 15492 24448 15556 24452
rect 18252 24508 18316 24512
rect 18252 24452 18256 24508
rect 18256 24452 18312 24508
rect 18312 24452 18316 24508
rect 18252 24448 18316 24452
rect 18332 24508 18396 24512
rect 18332 24452 18336 24508
rect 18336 24452 18392 24508
rect 18392 24452 18396 24508
rect 18332 24448 18396 24452
rect 18412 24508 18476 24512
rect 18412 24452 18416 24508
rect 18416 24452 18472 24508
rect 18472 24452 18476 24508
rect 18412 24448 18476 24452
rect 18492 24508 18556 24512
rect 18492 24452 18496 24508
rect 18496 24452 18552 24508
rect 18552 24452 18556 24508
rect 18492 24448 18556 24452
rect 21252 24508 21316 24512
rect 21252 24452 21256 24508
rect 21256 24452 21312 24508
rect 21312 24452 21316 24508
rect 21252 24448 21316 24452
rect 21332 24508 21396 24512
rect 21332 24452 21336 24508
rect 21336 24452 21392 24508
rect 21392 24452 21396 24508
rect 21332 24448 21396 24452
rect 21412 24508 21476 24512
rect 21412 24452 21416 24508
rect 21416 24452 21472 24508
rect 21472 24452 21476 24508
rect 21412 24448 21476 24452
rect 21492 24508 21556 24512
rect 21492 24452 21496 24508
rect 21496 24452 21552 24508
rect 21552 24452 21556 24508
rect 21492 24448 21556 24452
rect 24252 24508 24316 24512
rect 24252 24452 24256 24508
rect 24256 24452 24312 24508
rect 24312 24452 24316 24508
rect 24252 24448 24316 24452
rect 24332 24508 24396 24512
rect 24332 24452 24336 24508
rect 24336 24452 24392 24508
rect 24392 24452 24396 24508
rect 24332 24448 24396 24452
rect 24412 24508 24476 24512
rect 24412 24452 24416 24508
rect 24416 24452 24472 24508
rect 24472 24452 24476 24508
rect 24412 24448 24476 24452
rect 24492 24508 24556 24512
rect 24492 24452 24496 24508
rect 24496 24452 24552 24508
rect 24552 24452 24556 24508
rect 24492 24448 24556 24452
rect 27252 24508 27316 24512
rect 27252 24452 27256 24508
rect 27256 24452 27312 24508
rect 27312 24452 27316 24508
rect 27252 24448 27316 24452
rect 27332 24508 27396 24512
rect 27332 24452 27336 24508
rect 27336 24452 27392 24508
rect 27392 24452 27396 24508
rect 27332 24448 27396 24452
rect 27412 24508 27476 24512
rect 27412 24452 27416 24508
rect 27416 24452 27472 24508
rect 27472 24452 27476 24508
rect 27412 24448 27476 24452
rect 27492 24508 27556 24512
rect 27492 24452 27496 24508
rect 27496 24452 27552 24508
rect 27552 24452 27556 24508
rect 27492 24448 27556 24452
rect 1752 23964 1816 23968
rect 1752 23908 1756 23964
rect 1756 23908 1812 23964
rect 1812 23908 1816 23964
rect 1752 23904 1816 23908
rect 1832 23964 1896 23968
rect 1832 23908 1836 23964
rect 1836 23908 1892 23964
rect 1892 23908 1896 23964
rect 1832 23904 1896 23908
rect 1912 23964 1976 23968
rect 1912 23908 1916 23964
rect 1916 23908 1972 23964
rect 1972 23908 1976 23964
rect 1912 23904 1976 23908
rect 1992 23964 2056 23968
rect 1992 23908 1996 23964
rect 1996 23908 2052 23964
rect 2052 23908 2056 23964
rect 1992 23904 2056 23908
rect 4752 23964 4816 23968
rect 4752 23908 4756 23964
rect 4756 23908 4812 23964
rect 4812 23908 4816 23964
rect 4752 23904 4816 23908
rect 4832 23964 4896 23968
rect 4832 23908 4836 23964
rect 4836 23908 4892 23964
rect 4892 23908 4896 23964
rect 4832 23904 4896 23908
rect 4912 23964 4976 23968
rect 4912 23908 4916 23964
rect 4916 23908 4972 23964
rect 4972 23908 4976 23964
rect 4912 23904 4976 23908
rect 4992 23964 5056 23968
rect 4992 23908 4996 23964
rect 4996 23908 5052 23964
rect 5052 23908 5056 23964
rect 4992 23904 5056 23908
rect 7752 23964 7816 23968
rect 7752 23908 7756 23964
rect 7756 23908 7812 23964
rect 7812 23908 7816 23964
rect 7752 23904 7816 23908
rect 7832 23964 7896 23968
rect 7832 23908 7836 23964
rect 7836 23908 7892 23964
rect 7892 23908 7896 23964
rect 7832 23904 7896 23908
rect 7912 23964 7976 23968
rect 7912 23908 7916 23964
rect 7916 23908 7972 23964
rect 7972 23908 7976 23964
rect 7912 23904 7976 23908
rect 7992 23964 8056 23968
rect 7992 23908 7996 23964
rect 7996 23908 8052 23964
rect 8052 23908 8056 23964
rect 7992 23904 8056 23908
rect 10752 23964 10816 23968
rect 10752 23908 10756 23964
rect 10756 23908 10812 23964
rect 10812 23908 10816 23964
rect 10752 23904 10816 23908
rect 10832 23964 10896 23968
rect 10832 23908 10836 23964
rect 10836 23908 10892 23964
rect 10892 23908 10896 23964
rect 10832 23904 10896 23908
rect 10912 23964 10976 23968
rect 10912 23908 10916 23964
rect 10916 23908 10972 23964
rect 10972 23908 10976 23964
rect 10912 23904 10976 23908
rect 10992 23964 11056 23968
rect 10992 23908 10996 23964
rect 10996 23908 11052 23964
rect 11052 23908 11056 23964
rect 10992 23904 11056 23908
rect 13752 23964 13816 23968
rect 13752 23908 13756 23964
rect 13756 23908 13812 23964
rect 13812 23908 13816 23964
rect 13752 23904 13816 23908
rect 13832 23964 13896 23968
rect 13832 23908 13836 23964
rect 13836 23908 13892 23964
rect 13892 23908 13896 23964
rect 13832 23904 13896 23908
rect 13912 23964 13976 23968
rect 13912 23908 13916 23964
rect 13916 23908 13972 23964
rect 13972 23908 13976 23964
rect 13912 23904 13976 23908
rect 13992 23964 14056 23968
rect 13992 23908 13996 23964
rect 13996 23908 14052 23964
rect 14052 23908 14056 23964
rect 13992 23904 14056 23908
rect 16752 23964 16816 23968
rect 16752 23908 16756 23964
rect 16756 23908 16812 23964
rect 16812 23908 16816 23964
rect 16752 23904 16816 23908
rect 16832 23964 16896 23968
rect 16832 23908 16836 23964
rect 16836 23908 16892 23964
rect 16892 23908 16896 23964
rect 16832 23904 16896 23908
rect 16912 23964 16976 23968
rect 16912 23908 16916 23964
rect 16916 23908 16972 23964
rect 16972 23908 16976 23964
rect 16912 23904 16976 23908
rect 16992 23964 17056 23968
rect 16992 23908 16996 23964
rect 16996 23908 17052 23964
rect 17052 23908 17056 23964
rect 16992 23904 17056 23908
rect 19752 23964 19816 23968
rect 19752 23908 19756 23964
rect 19756 23908 19812 23964
rect 19812 23908 19816 23964
rect 19752 23904 19816 23908
rect 19832 23964 19896 23968
rect 19832 23908 19836 23964
rect 19836 23908 19892 23964
rect 19892 23908 19896 23964
rect 19832 23904 19896 23908
rect 19912 23964 19976 23968
rect 19912 23908 19916 23964
rect 19916 23908 19972 23964
rect 19972 23908 19976 23964
rect 19912 23904 19976 23908
rect 19992 23964 20056 23968
rect 19992 23908 19996 23964
rect 19996 23908 20052 23964
rect 20052 23908 20056 23964
rect 19992 23904 20056 23908
rect 22752 23964 22816 23968
rect 22752 23908 22756 23964
rect 22756 23908 22812 23964
rect 22812 23908 22816 23964
rect 22752 23904 22816 23908
rect 22832 23964 22896 23968
rect 22832 23908 22836 23964
rect 22836 23908 22892 23964
rect 22892 23908 22896 23964
rect 22832 23904 22896 23908
rect 22912 23964 22976 23968
rect 22912 23908 22916 23964
rect 22916 23908 22972 23964
rect 22972 23908 22976 23964
rect 22912 23904 22976 23908
rect 22992 23964 23056 23968
rect 22992 23908 22996 23964
rect 22996 23908 23052 23964
rect 23052 23908 23056 23964
rect 22992 23904 23056 23908
rect 25752 23964 25816 23968
rect 25752 23908 25756 23964
rect 25756 23908 25812 23964
rect 25812 23908 25816 23964
rect 25752 23904 25816 23908
rect 25832 23964 25896 23968
rect 25832 23908 25836 23964
rect 25836 23908 25892 23964
rect 25892 23908 25896 23964
rect 25832 23904 25896 23908
rect 25912 23964 25976 23968
rect 25912 23908 25916 23964
rect 25916 23908 25972 23964
rect 25972 23908 25976 23964
rect 25912 23904 25976 23908
rect 25992 23964 26056 23968
rect 25992 23908 25996 23964
rect 25996 23908 26052 23964
rect 26052 23908 26056 23964
rect 25992 23904 26056 23908
rect 3252 23420 3316 23424
rect 3252 23364 3256 23420
rect 3256 23364 3312 23420
rect 3312 23364 3316 23420
rect 3252 23360 3316 23364
rect 3332 23420 3396 23424
rect 3332 23364 3336 23420
rect 3336 23364 3392 23420
rect 3392 23364 3396 23420
rect 3332 23360 3396 23364
rect 3412 23420 3476 23424
rect 3412 23364 3416 23420
rect 3416 23364 3472 23420
rect 3472 23364 3476 23420
rect 3412 23360 3476 23364
rect 3492 23420 3556 23424
rect 3492 23364 3496 23420
rect 3496 23364 3552 23420
rect 3552 23364 3556 23420
rect 3492 23360 3556 23364
rect 6252 23420 6316 23424
rect 6252 23364 6256 23420
rect 6256 23364 6312 23420
rect 6312 23364 6316 23420
rect 6252 23360 6316 23364
rect 6332 23420 6396 23424
rect 6332 23364 6336 23420
rect 6336 23364 6392 23420
rect 6392 23364 6396 23420
rect 6332 23360 6396 23364
rect 6412 23420 6476 23424
rect 6412 23364 6416 23420
rect 6416 23364 6472 23420
rect 6472 23364 6476 23420
rect 6412 23360 6476 23364
rect 6492 23420 6556 23424
rect 6492 23364 6496 23420
rect 6496 23364 6552 23420
rect 6552 23364 6556 23420
rect 6492 23360 6556 23364
rect 9252 23420 9316 23424
rect 9252 23364 9256 23420
rect 9256 23364 9312 23420
rect 9312 23364 9316 23420
rect 9252 23360 9316 23364
rect 9332 23420 9396 23424
rect 9332 23364 9336 23420
rect 9336 23364 9392 23420
rect 9392 23364 9396 23420
rect 9332 23360 9396 23364
rect 9412 23420 9476 23424
rect 9412 23364 9416 23420
rect 9416 23364 9472 23420
rect 9472 23364 9476 23420
rect 9412 23360 9476 23364
rect 9492 23420 9556 23424
rect 9492 23364 9496 23420
rect 9496 23364 9552 23420
rect 9552 23364 9556 23420
rect 9492 23360 9556 23364
rect 12252 23420 12316 23424
rect 12252 23364 12256 23420
rect 12256 23364 12312 23420
rect 12312 23364 12316 23420
rect 12252 23360 12316 23364
rect 12332 23420 12396 23424
rect 12332 23364 12336 23420
rect 12336 23364 12392 23420
rect 12392 23364 12396 23420
rect 12332 23360 12396 23364
rect 12412 23420 12476 23424
rect 12412 23364 12416 23420
rect 12416 23364 12472 23420
rect 12472 23364 12476 23420
rect 12412 23360 12476 23364
rect 12492 23420 12556 23424
rect 12492 23364 12496 23420
rect 12496 23364 12552 23420
rect 12552 23364 12556 23420
rect 12492 23360 12556 23364
rect 15252 23420 15316 23424
rect 15252 23364 15256 23420
rect 15256 23364 15312 23420
rect 15312 23364 15316 23420
rect 15252 23360 15316 23364
rect 15332 23420 15396 23424
rect 15332 23364 15336 23420
rect 15336 23364 15392 23420
rect 15392 23364 15396 23420
rect 15332 23360 15396 23364
rect 15412 23420 15476 23424
rect 15412 23364 15416 23420
rect 15416 23364 15472 23420
rect 15472 23364 15476 23420
rect 15412 23360 15476 23364
rect 15492 23420 15556 23424
rect 15492 23364 15496 23420
rect 15496 23364 15552 23420
rect 15552 23364 15556 23420
rect 15492 23360 15556 23364
rect 18252 23420 18316 23424
rect 18252 23364 18256 23420
rect 18256 23364 18312 23420
rect 18312 23364 18316 23420
rect 18252 23360 18316 23364
rect 18332 23420 18396 23424
rect 18332 23364 18336 23420
rect 18336 23364 18392 23420
rect 18392 23364 18396 23420
rect 18332 23360 18396 23364
rect 18412 23420 18476 23424
rect 18412 23364 18416 23420
rect 18416 23364 18472 23420
rect 18472 23364 18476 23420
rect 18412 23360 18476 23364
rect 18492 23420 18556 23424
rect 18492 23364 18496 23420
rect 18496 23364 18552 23420
rect 18552 23364 18556 23420
rect 18492 23360 18556 23364
rect 21252 23420 21316 23424
rect 21252 23364 21256 23420
rect 21256 23364 21312 23420
rect 21312 23364 21316 23420
rect 21252 23360 21316 23364
rect 21332 23420 21396 23424
rect 21332 23364 21336 23420
rect 21336 23364 21392 23420
rect 21392 23364 21396 23420
rect 21332 23360 21396 23364
rect 21412 23420 21476 23424
rect 21412 23364 21416 23420
rect 21416 23364 21472 23420
rect 21472 23364 21476 23420
rect 21412 23360 21476 23364
rect 21492 23420 21556 23424
rect 21492 23364 21496 23420
rect 21496 23364 21552 23420
rect 21552 23364 21556 23420
rect 21492 23360 21556 23364
rect 24252 23420 24316 23424
rect 24252 23364 24256 23420
rect 24256 23364 24312 23420
rect 24312 23364 24316 23420
rect 24252 23360 24316 23364
rect 24332 23420 24396 23424
rect 24332 23364 24336 23420
rect 24336 23364 24392 23420
rect 24392 23364 24396 23420
rect 24332 23360 24396 23364
rect 24412 23420 24476 23424
rect 24412 23364 24416 23420
rect 24416 23364 24472 23420
rect 24472 23364 24476 23420
rect 24412 23360 24476 23364
rect 24492 23420 24556 23424
rect 24492 23364 24496 23420
rect 24496 23364 24552 23420
rect 24552 23364 24556 23420
rect 24492 23360 24556 23364
rect 27252 23420 27316 23424
rect 27252 23364 27256 23420
rect 27256 23364 27312 23420
rect 27312 23364 27316 23420
rect 27252 23360 27316 23364
rect 27332 23420 27396 23424
rect 27332 23364 27336 23420
rect 27336 23364 27392 23420
rect 27392 23364 27396 23420
rect 27332 23360 27396 23364
rect 27412 23420 27476 23424
rect 27412 23364 27416 23420
rect 27416 23364 27472 23420
rect 27472 23364 27476 23420
rect 27412 23360 27476 23364
rect 27492 23420 27556 23424
rect 27492 23364 27496 23420
rect 27496 23364 27552 23420
rect 27552 23364 27556 23420
rect 27492 23360 27556 23364
rect 1752 22876 1816 22880
rect 1752 22820 1756 22876
rect 1756 22820 1812 22876
rect 1812 22820 1816 22876
rect 1752 22816 1816 22820
rect 1832 22876 1896 22880
rect 1832 22820 1836 22876
rect 1836 22820 1892 22876
rect 1892 22820 1896 22876
rect 1832 22816 1896 22820
rect 1912 22876 1976 22880
rect 1912 22820 1916 22876
rect 1916 22820 1972 22876
rect 1972 22820 1976 22876
rect 1912 22816 1976 22820
rect 1992 22876 2056 22880
rect 1992 22820 1996 22876
rect 1996 22820 2052 22876
rect 2052 22820 2056 22876
rect 1992 22816 2056 22820
rect 4752 22876 4816 22880
rect 4752 22820 4756 22876
rect 4756 22820 4812 22876
rect 4812 22820 4816 22876
rect 4752 22816 4816 22820
rect 4832 22876 4896 22880
rect 4832 22820 4836 22876
rect 4836 22820 4892 22876
rect 4892 22820 4896 22876
rect 4832 22816 4896 22820
rect 4912 22876 4976 22880
rect 4912 22820 4916 22876
rect 4916 22820 4972 22876
rect 4972 22820 4976 22876
rect 4912 22816 4976 22820
rect 4992 22876 5056 22880
rect 4992 22820 4996 22876
rect 4996 22820 5052 22876
rect 5052 22820 5056 22876
rect 4992 22816 5056 22820
rect 7752 22876 7816 22880
rect 7752 22820 7756 22876
rect 7756 22820 7812 22876
rect 7812 22820 7816 22876
rect 7752 22816 7816 22820
rect 7832 22876 7896 22880
rect 7832 22820 7836 22876
rect 7836 22820 7892 22876
rect 7892 22820 7896 22876
rect 7832 22816 7896 22820
rect 7912 22876 7976 22880
rect 7912 22820 7916 22876
rect 7916 22820 7972 22876
rect 7972 22820 7976 22876
rect 7912 22816 7976 22820
rect 7992 22876 8056 22880
rect 7992 22820 7996 22876
rect 7996 22820 8052 22876
rect 8052 22820 8056 22876
rect 7992 22816 8056 22820
rect 10752 22876 10816 22880
rect 10752 22820 10756 22876
rect 10756 22820 10812 22876
rect 10812 22820 10816 22876
rect 10752 22816 10816 22820
rect 10832 22876 10896 22880
rect 10832 22820 10836 22876
rect 10836 22820 10892 22876
rect 10892 22820 10896 22876
rect 10832 22816 10896 22820
rect 10912 22876 10976 22880
rect 10912 22820 10916 22876
rect 10916 22820 10972 22876
rect 10972 22820 10976 22876
rect 10912 22816 10976 22820
rect 10992 22876 11056 22880
rect 10992 22820 10996 22876
rect 10996 22820 11052 22876
rect 11052 22820 11056 22876
rect 10992 22816 11056 22820
rect 13752 22876 13816 22880
rect 13752 22820 13756 22876
rect 13756 22820 13812 22876
rect 13812 22820 13816 22876
rect 13752 22816 13816 22820
rect 13832 22876 13896 22880
rect 13832 22820 13836 22876
rect 13836 22820 13892 22876
rect 13892 22820 13896 22876
rect 13832 22816 13896 22820
rect 13912 22876 13976 22880
rect 13912 22820 13916 22876
rect 13916 22820 13972 22876
rect 13972 22820 13976 22876
rect 13912 22816 13976 22820
rect 13992 22876 14056 22880
rect 13992 22820 13996 22876
rect 13996 22820 14052 22876
rect 14052 22820 14056 22876
rect 13992 22816 14056 22820
rect 16752 22876 16816 22880
rect 16752 22820 16756 22876
rect 16756 22820 16812 22876
rect 16812 22820 16816 22876
rect 16752 22816 16816 22820
rect 16832 22876 16896 22880
rect 16832 22820 16836 22876
rect 16836 22820 16892 22876
rect 16892 22820 16896 22876
rect 16832 22816 16896 22820
rect 16912 22876 16976 22880
rect 16912 22820 16916 22876
rect 16916 22820 16972 22876
rect 16972 22820 16976 22876
rect 16912 22816 16976 22820
rect 16992 22876 17056 22880
rect 16992 22820 16996 22876
rect 16996 22820 17052 22876
rect 17052 22820 17056 22876
rect 16992 22816 17056 22820
rect 19752 22876 19816 22880
rect 19752 22820 19756 22876
rect 19756 22820 19812 22876
rect 19812 22820 19816 22876
rect 19752 22816 19816 22820
rect 19832 22876 19896 22880
rect 19832 22820 19836 22876
rect 19836 22820 19892 22876
rect 19892 22820 19896 22876
rect 19832 22816 19896 22820
rect 19912 22876 19976 22880
rect 19912 22820 19916 22876
rect 19916 22820 19972 22876
rect 19972 22820 19976 22876
rect 19912 22816 19976 22820
rect 19992 22876 20056 22880
rect 19992 22820 19996 22876
rect 19996 22820 20052 22876
rect 20052 22820 20056 22876
rect 19992 22816 20056 22820
rect 22752 22876 22816 22880
rect 22752 22820 22756 22876
rect 22756 22820 22812 22876
rect 22812 22820 22816 22876
rect 22752 22816 22816 22820
rect 22832 22876 22896 22880
rect 22832 22820 22836 22876
rect 22836 22820 22892 22876
rect 22892 22820 22896 22876
rect 22832 22816 22896 22820
rect 22912 22876 22976 22880
rect 22912 22820 22916 22876
rect 22916 22820 22972 22876
rect 22972 22820 22976 22876
rect 22912 22816 22976 22820
rect 22992 22876 23056 22880
rect 22992 22820 22996 22876
rect 22996 22820 23052 22876
rect 23052 22820 23056 22876
rect 22992 22816 23056 22820
rect 25752 22876 25816 22880
rect 25752 22820 25756 22876
rect 25756 22820 25812 22876
rect 25812 22820 25816 22876
rect 25752 22816 25816 22820
rect 25832 22876 25896 22880
rect 25832 22820 25836 22876
rect 25836 22820 25892 22876
rect 25892 22820 25896 22876
rect 25832 22816 25896 22820
rect 25912 22876 25976 22880
rect 25912 22820 25916 22876
rect 25916 22820 25972 22876
rect 25972 22820 25976 22876
rect 25912 22816 25976 22820
rect 25992 22876 26056 22880
rect 25992 22820 25996 22876
rect 25996 22820 26052 22876
rect 26052 22820 26056 22876
rect 25992 22816 26056 22820
rect 3252 22332 3316 22336
rect 3252 22276 3256 22332
rect 3256 22276 3312 22332
rect 3312 22276 3316 22332
rect 3252 22272 3316 22276
rect 3332 22332 3396 22336
rect 3332 22276 3336 22332
rect 3336 22276 3392 22332
rect 3392 22276 3396 22332
rect 3332 22272 3396 22276
rect 3412 22332 3476 22336
rect 3412 22276 3416 22332
rect 3416 22276 3472 22332
rect 3472 22276 3476 22332
rect 3412 22272 3476 22276
rect 3492 22332 3556 22336
rect 3492 22276 3496 22332
rect 3496 22276 3552 22332
rect 3552 22276 3556 22332
rect 3492 22272 3556 22276
rect 6252 22332 6316 22336
rect 6252 22276 6256 22332
rect 6256 22276 6312 22332
rect 6312 22276 6316 22332
rect 6252 22272 6316 22276
rect 6332 22332 6396 22336
rect 6332 22276 6336 22332
rect 6336 22276 6392 22332
rect 6392 22276 6396 22332
rect 6332 22272 6396 22276
rect 6412 22332 6476 22336
rect 6412 22276 6416 22332
rect 6416 22276 6472 22332
rect 6472 22276 6476 22332
rect 6412 22272 6476 22276
rect 6492 22332 6556 22336
rect 6492 22276 6496 22332
rect 6496 22276 6552 22332
rect 6552 22276 6556 22332
rect 6492 22272 6556 22276
rect 9252 22332 9316 22336
rect 9252 22276 9256 22332
rect 9256 22276 9312 22332
rect 9312 22276 9316 22332
rect 9252 22272 9316 22276
rect 9332 22332 9396 22336
rect 9332 22276 9336 22332
rect 9336 22276 9392 22332
rect 9392 22276 9396 22332
rect 9332 22272 9396 22276
rect 9412 22332 9476 22336
rect 9412 22276 9416 22332
rect 9416 22276 9472 22332
rect 9472 22276 9476 22332
rect 9412 22272 9476 22276
rect 9492 22332 9556 22336
rect 9492 22276 9496 22332
rect 9496 22276 9552 22332
rect 9552 22276 9556 22332
rect 9492 22272 9556 22276
rect 12252 22332 12316 22336
rect 12252 22276 12256 22332
rect 12256 22276 12312 22332
rect 12312 22276 12316 22332
rect 12252 22272 12316 22276
rect 12332 22332 12396 22336
rect 12332 22276 12336 22332
rect 12336 22276 12392 22332
rect 12392 22276 12396 22332
rect 12332 22272 12396 22276
rect 12412 22332 12476 22336
rect 12412 22276 12416 22332
rect 12416 22276 12472 22332
rect 12472 22276 12476 22332
rect 12412 22272 12476 22276
rect 12492 22332 12556 22336
rect 12492 22276 12496 22332
rect 12496 22276 12552 22332
rect 12552 22276 12556 22332
rect 12492 22272 12556 22276
rect 15252 22332 15316 22336
rect 15252 22276 15256 22332
rect 15256 22276 15312 22332
rect 15312 22276 15316 22332
rect 15252 22272 15316 22276
rect 15332 22332 15396 22336
rect 15332 22276 15336 22332
rect 15336 22276 15392 22332
rect 15392 22276 15396 22332
rect 15332 22272 15396 22276
rect 15412 22332 15476 22336
rect 15412 22276 15416 22332
rect 15416 22276 15472 22332
rect 15472 22276 15476 22332
rect 15412 22272 15476 22276
rect 15492 22332 15556 22336
rect 15492 22276 15496 22332
rect 15496 22276 15552 22332
rect 15552 22276 15556 22332
rect 15492 22272 15556 22276
rect 18252 22332 18316 22336
rect 18252 22276 18256 22332
rect 18256 22276 18312 22332
rect 18312 22276 18316 22332
rect 18252 22272 18316 22276
rect 18332 22332 18396 22336
rect 18332 22276 18336 22332
rect 18336 22276 18392 22332
rect 18392 22276 18396 22332
rect 18332 22272 18396 22276
rect 18412 22332 18476 22336
rect 18412 22276 18416 22332
rect 18416 22276 18472 22332
rect 18472 22276 18476 22332
rect 18412 22272 18476 22276
rect 18492 22332 18556 22336
rect 18492 22276 18496 22332
rect 18496 22276 18552 22332
rect 18552 22276 18556 22332
rect 18492 22272 18556 22276
rect 21252 22332 21316 22336
rect 21252 22276 21256 22332
rect 21256 22276 21312 22332
rect 21312 22276 21316 22332
rect 21252 22272 21316 22276
rect 21332 22332 21396 22336
rect 21332 22276 21336 22332
rect 21336 22276 21392 22332
rect 21392 22276 21396 22332
rect 21332 22272 21396 22276
rect 21412 22332 21476 22336
rect 21412 22276 21416 22332
rect 21416 22276 21472 22332
rect 21472 22276 21476 22332
rect 21412 22272 21476 22276
rect 21492 22332 21556 22336
rect 21492 22276 21496 22332
rect 21496 22276 21552 22332
rect 21552 22276 21556 22332
rect 21492 22272 21556 22276
rect 24252 22332 24316 22336
rect 24252 22276 24256 22332
rect 24256 22276 24312 22332
rect 24312 22276 24316 22332
rect 24252 22272 24316 22276
rect 24332 22332 24396 22336
rect 24332 22276 24336 22332
rect 24336 22276 24392 22332
rect 24392 22276 24396 22332
rect 24332 22272 24396 22276
rect 24412 22332 24476 22336
rect 24412 22276 24416 22332
rect 24416 22276 24472 22332
rect 24472 22276 24476 22332
rect 24412 22272 24476 22276
rect 24492 22332 24556 22336
rect 24492 22276 24496 22332
rect 24496 22276 24552 22332
rect 24552 22276 24556 22332
rect 24492 22272 24556 22276
rect 27252 22332 27316 22336
rect 27252 22276 27256 22332
rect 27256 22276 27312 22332
rect 27312 22276 27316 22332
rect 27252 22272 27316 22276
rect 27332 22332 27396 22336
rect 27332 22276 27336 22332
rect 27336 22276 27392 22332
rect 27392 22276 27396 22332
rect 27332 22272 27396 22276
rect 27412 22332 27476 22336
rect 27412 22276 27416 22332
rect 27416 22276 27472 22332
rect 27472 22276 27476 22332
rect 27412 22272 27476 22276
rect 27492 22332 27556 22336
rect 27492 22276 27496 22332
rect 27496 22276 27552 22332
rect 27552 22276 27556 22332
rect 27492 22272 27556 22276
rect 1752 21788 1816 21792
rect 1752 21732 1756 21788
rect 1756 21732 1812 21788
rect 1812 21732 1816 21788
rect 1752 21728 1816 21732
rect 1832 21788 1896 21792
rect 1832 21732 1836 21788
rect 1836 21732 1892 21788
rect 1892 21732 1896 21788
rect 1832 21728 1896 21732
rect 1912 21788 1976 21792
rect 1912 21732 1916 21788
rect 1916 21732 1972 21788
rect 1972 21732 1976 21788
rect 1912 21728 1976 21732
rect 1992 21788 2056 21792
rect 1992 21732 1996 21788
rect 1996 21732 2052 21788
rect 2052 21732 2056 21788
rect 1992 21728 2056 21732
rect 4752 21788 4816 21792
rect 4752 21732 4756 21788
rect 4756 21732 4812 21788
rect 4812 21732 4816 21788
rect 4752 21728 4816 21732
rect 4832 21788 4896 21792
rect 4832 21732 4836 21788
rect 4836 21732 4892 21788
rect 4892 21732 4896 21788
rect 4832 21728 4896 21732
rect 4912 21788 4976 21792
rect 4912 21732 4916 21788
rect 4916 21732 4972 21788
rect 4972 21732 4976 21788
rect 4912 21728 4976 21732
rect 4992 21788 5056 21792
rect 4992 21732 4996 21788
rect 4996 21732 5052 21788
rect 5052 21732 5056 21788
rect 4992 21728 5056 21732
rect 7752 21788 7816 21792
rect 7752 21732 7756 21788
rect 7756 21732 7812 21788
rect 7812 21732 7816 21788
rect 7752 21728 7816 21732
rect 7832 21788 7896 21792
rect 7832 21732 7836 21788
rect 7836 21732 7892 21788
rect 7892 21732 7896 21788
rect 7832 21728 7896 21732
rect 7912 21788 7976 21792
rect 7912 21732 7916 21788
rect 7916 21732 7972 21788
rect 7972 21732 7976 21788
rect 7912 21728 7976 21732
rect 7992 21788 8056 21792
rect 7992 21732 7996 21788
rect 7996 21732 8052 21788
rect 8052 21732 8056 21788
rect 7992 21728 8056 21732
rect 10752 21788 10816 21792
rect 10752 21732 10756 21788
rect 10756 21732 10812 21788
rect 10812 21732 10816 21788
rect 10752 21728 10816 21732
rect 10832 21788 10896 21792
rect 10832 21732 10836 21788
rect 10836 21732 10892 21788
rect 10892 21732 10896 21788
rect 10832 21728 10896 21732
rect 10912 21788 10976 21792
rect 10912 21732 10916 21788
rect 10916 21732 10972 21788
rect 10972 21732 10976 21788
rect 10912 21728 10976 21732
rect 10992 21788 11056 21792
rect 10992 21732 10996 21788
rect 10996 21732 11052 21788
rect 11052 21732 11056 21788
rect 10992 21728 11056 21732
rect 13752 21788 13816 21792
rect 13752 21732 13756 21788
rect 13756 21732 13812 21788
rect 13812 21732 13816 21788
rect 13752 21728 13816 21732
rect 13832 21788 13896 21792
rect 13832 21732 13836 21788
rect 13836 21732 13892 21788
rect 13892 21732 13896 21788
rect 13832 21728 13896 21732
rect 13912 21788 13976 21792
rect 13912 21732 13916 21788
rect 13916 21732 13972 21788
rect 13972 21732 13976 21788
rect 13912 21728 13976 21732
rect 13992 21788 14056 21792
rect 13992 21732 13996 21788
rect 13996 21732 14052 21788
rect 14052 21732 14056 21788
rect 13992 21728 14056 21732
rect 16752 21788 16816 21792
rect 16752 21732 16756 21788
rect 16756 21732 16812 21788
rect 16812 21732 16816 21788
rect 16752 21728 16816 21732
rect 16832 21788 16896 21792
rect 16832 21732 16836 21788
rect 16836 21732 16892 21788
rect 16892 21732 16896 21788
rect 16832 21728 16896 21732
rect 16912 21788 16976 21792
rect 16912 21732 16916 21788
rect 16916 21732 16972 21788
rect 16972 21732 16976 21788
rect 16912 21728 16976 21732
rect 16992 21788 17056 21792
rect 16992 21732 16996 21788
rect 16996 21732 17052 21788
rect 17052 21732 17056 21788
rect 16992 21728 17056 21732
rect 19752 21788 19816 21792
rect 19752 21732 19756 21788
rect 19756 21732 19812 21788
rect 19812 21732 19816 21788
rect 19752 21728 19816 21732
rect 19832 21788 19896 21792
rect 19832 21732 19836 21788
rect 19836 21732 19892 21788
rect 19892 21732 19896 21788
rect 19832 21728 19896 21732
rect 19912 21788 19976 21792
rect 19912 21732 19916 21788
rect 19916 21732 19972 21788
rect 19972 21732 19976 21788
rect 19912 21728 19976 21732
rect 19992 21788 20056 21792
rect 19992 21732 19996 21788
rect 19996 21732 20052 21788
rect 20052 21732 20056 21788
rect 19992 21728 20056 21732
rect 22752 21788 22816 21792
rect 22752 21732 22756 21788
rect 22756 21732 22812 21788
rect 22812 21732 22816 21788
rect 22752 21728 22816 21732
rect 22832 21788 22896 21792
rect 22832 21732 22836 21788
rect 22836 21732 22892 21788
rect 22892 21732 22896 21788
rect 22832 21728 22896 21732
rect 22912 21788 22976 21792
rect 22912 21732 22916 21788
rect 22916 21732 22972 21788
rect 22972 21732 22976 21788
rect 22912 21728 22976 21732
rect 22992 21788 23056 21792
rect 22992 21732 22996 21788
rect 22996 21732 23052 21788
rect 23052 21732 23056 21788
rect 22992 21728 23056 21732
rect 25752 21788 25816 21792
rect 25752 21732 25756 21788
rect 25756 21732 25812 21788
rect 25812 21732 25816 21788
rect 25752 21728 25816 21732
rect 25832 21788 25896 21792
rect 25832 21732 25836 21788
rect 25836 21732 25892 21788
rect 25892 21732 25896 21788
rect 25832 21728 25896 21732
rect 25912 21788 25976 21792
rect 25912 21732 25916 21788
rect 25916 21732 25972 21788
rect 25972 21732 25976 21788
rect 25912 21728 25976 21732
rect 25992 21788 26056 21792
rect 25992 21732 25996 21788
rect 25996 21732 26052 21788
rect 26052 21732 26056 21788
rect 25992 21728 26056 21732
rect 3252 21244 3316 21248
rect 3252 21188 3256 21244
rect 3256 21188 3312 21244
rect 3312 21188 3316 21244
rect 3252 21184 3316 21188
rect 3332 21244 3396 21248
rect 3332 21188 3336 21244
rect 3336 21188 3392 21244
rect 3392 21188 3396 21244
rect 3332 21184 3396 21188
rect 3412 21244 3476 21248
rect 3412 21188 3416 21244
rect 3416 21188 3472 21244
rect 3472 21188 3476 21244
rect 3412 21184 3476 21188
rect 3492 21244 3556 21248
rect 3492 21188 3496 21244
rect 3496 21188 3552 21244
rect 3552 21188 3556 21244
rect 3492 21184 3556 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 6412 21244 6476 21248
rect 6412 21188 6416 21244
rect 6416 21188 6472 21244
rect 6472 21188 6476 21244
rect 6412 21184 6476 21188
rect 6492 21244 6556 21248
rect 6492 21188 6496 21244
rect 6496 21188 6552 21244
rect 6552 21188 6556 21244
rect 6492 21184 6556 21188
rect 9252 21244 9316 21248
rect 9252 21188 9256 21244
rect 9256 21188 9312 21244
rect 9312 21188 9316 21244
rect 9252 21184 9316 21188
rect 9332 21244 9396 21248
rect 9332 21188 9336 21244
rect 9336 21188 9392 21244
rect 9392 21188 9396 21244
rect 9332 21184 9396 21188
rect 9412 21244 9476 21248
rect 9412 21188 9416 21244
rect 9416 21188 9472 21244
rect 9472 21188 9476 21244
rect 9412 21184 9476 21188
rect 9492 21244 9556 21248
rect 9492 21188 9496 21244
rect 9496 21188 9552 21244
rect 9552 21188 9556 21244
rect 9492 21184 9556 21188
rect 12252 21244 12316 21248
rect 12252 21188 12256 21244
rect 12256 21188 12312 21244
rect 12312 21188 12316 21244
rect 12252 21184 12316 21188
rect 12332 21244 12396 21248
rect 12332 21188 12336 21244
rect 12336 21188 12392 21244
rect 12392 21188 12396 21244
rect 12332 21184 12396 21188
rect 12412 21244 12476 21248
rect 12412 21188 12416 21244
rect 12416 21188 12472 21244
rect 12472 21188 12476 21244
rect 12412 21184 12476 21188
rect 12492 21244 12556 21248
rect 12492 21188 12496 21244
rect 12496 21188 12552 21244
rect 12552 21188 12556 21244
rect 12492 21184 12556 21188
rect 15252 21244 15316 21248
rect 15252 21188 15256 21244
rect 15256 21188 15312 21244
rect 15312 21188 15316 21244
rect 15252 21184 15316 21188
rect 15332 21244 15396 21248
rect 15332 21188 15336 21244
rect 15336 21188 15392 21244
rect 15392 21188 15396 21244
rect 15332 21184 15396 21188
rect 15412 21244 15476 21248
rect 15412 21188 15416 21244
rect 15416 21188 15472 21244
rect 15472 21188 15476 21244
rect 15412 21184 15476 21188
rect 15492 21244 15556 21248
rect 15492 21188 15496 21244
rect 15496 21188 15552 21244
rect 15552 21188 15556 21244
rect 15492 21184 15556 21188
rect 18252 21244 18316 21248
rect 18252 21188 18256 21244
rect 18256 21188 18312 21244
rect 18312 21188 18316 21244
rect 18252 21184 18316 21188
rect 18332 21244 18396 21248
rect 18332 21188 18336 21244
rect 18336 21188 18392 21244
rect 18392 21188 18396 21244
rect 18332 21184 18396 21188
rect 18412 21244 18476 21248
rect 18412 21188 18416 21244
rect 18416 21188 18472 21244
rect 18472 21188 18476 21244
rect 18412 21184 18476 21188
rect 18492 21244 18556 21248
rect 18492 21188 18496 21244
rect 18496 21188 18552 21244
rect 18552 21188 18556 21244
rect 18492 21184 18556 21188
rect 21252 21244 21316 21248
rect 21252 21188 21256 21244
rect 21256 21188 21312 21244
rect 21312 21188 21316 21244
rect 21252 21184 21316 21188
rect 21332 21244 21396 21248
rect 21332 21188 21336 21244
rect 21336 21188 21392 21244
rect 21392 21188 21396 21244
rect 21332 21184 21396 21188
rect 21412 21244 21476 21248
rect 21412 21188 21416 21244
rect 21416 21188 21472 21244
rect 21472 21188 21476 21244
rect 21412 21184 21476 21188
rect 21492 21244 21556 21248
rect 21492 21188 21496 21244
rect 21496 21188 21552 21244
rect 21552 21188 21556 21244
rect 21492 21184 21556 21188
rect 24252 21244 24316 21248
rect 24252 21188 24256 21244
rect 24256 21188 24312 21244
rect 24312 21188 24316 21244
rect 24252 21184 24316 21188
rect 24332 21244 24396 21248
rect 24332 21188 24336 21244
rect 24336 21188 24392 21244
rect 24392 21188 24396 21244
rect 24332 21184 24396 21188
rect 24412 21244 24476 21248
rect 24412 21188 24416 21244
rect 24416 21188 24472 21244
rect 24472 21188 24476 21244
rect 24412 21184 24476 21188
rect 24492 21244 24556 21248
rect 24492 21188 24496 21244
rect 24496 21188 24552 21244
rect 24552 21188 24556 21244
rect 24492 21184 24556 21188
rect 27252 21244 27316 21248
rect 27252 21188 27256 21244
rect 27256 21188 27312 21244
rect 27312 21188 27316 21244
rect 27252 21184 27316 21188
rect 27332 21244 27396 21248
rect 27332 21188 27336 21244
rect 27336 21188 27392 21244
rect 27392 21188 27396 21244
rect 27332 21184 27396 21188
rect 27412 21244 27476 21248
rect 27412 21188 27416 21244
rect 27416 21188 27472 21244
rect 27472 21188 27476 21244
rect 27412 21184 27476 21188
rect 27492 21244 27556 21248
rect 27492 21188 27496 21244
rect 27496 21188 27552 21244
rect 27552 21188 27556 21244
rect 27492 21184 27556 21188
rect 1752 20700 1816 20704
rect 1752 20644 1756 20700
rect 1756 20644 1812 20700
rect 1812 20644 1816 20700
rect 1752 20640 1816 20644
rect 1832 20700 1896 20704
rect 1832 20644 1836 20700
rect 1836 20644 1892 20700
rect 1892 20644 1896 20700
rect 1832 20640 1896 20644
rect 1912 20700 1976 20704
rect 1912 20644 1916 20700
rect 1916 20644 1972 20700
rect 1972 20644 1976 20700
rect 1912 20640 1976 20644
rect 1992 20700 2056 20704
rect 1992 20644 1996 20700
rect 1996 20644 2052 20700
rect 2052 20644 2056 20700
rect 1992 20640 2056 20644
rect 4752 20700 4816 20704
rect 4752 20644 4756 20700
rect 4756 20644 4812 20700
rect 4812 20644 4816 20700
rect 4752 20640 4816 20644
rect 4832 20700 4896 20704
rect 4832 20644 4836 20700
rect 4836 20644 4892 20700
rect 4892 20644 4896 20700
rect 4832 20640 4896 20644
rect 4912 20700 4976 20704
rect 4912 20644 4916 20700
rect 4916 20644 4972 20700
rect 4972 20644 4976 20700
rect 4912 20640 4976 20644
rect 4992 20700 5056 20704
rect 4992 20644 4996 20700
rect 4996 20644 5052 20700
rect 5052 20644 5056 20700
rect 4992 20640 5056 20644
rect 7752 20700 7816 20704
rect 7752 20644 7756 20700
rect 7756 20644 7812 20700
rect 7812 20644 7816 20700
rect 7752 20640 7816 20644
rect 7832 20700 7896 20704
rect 7832 20644 7836 20700
rect 7836 20644 7892 20700
rect 7892 20644 7896 20700
rect 7832 20640 7896 20644
rect 7912 20700 7976 20704
rect 7912 20644 7916 20700
rect 7916 20644 7972 20700
rect 7972 20644 7976 20700
rect 7912 20640 7976 20644
rect 7992 20700 8056 20704
rect 7992 20644 7996 20700
rect 7996 20644 8052 20700
rect 8052 20644 8056 20700
rect 7992 20640 8056 20644
rect 10752 20700 10816 20704
rect 10752 20644 10756 20700
rect 10756 20644 10812 20700
rect 10812 20644 10816 20700
rect 10752 20640 10816 20644
rect 10832 20700 10896 20704
rect 10832 20644 10836 20700
rect 10836 20644 10892 20700
rect 10892 20644 10896 20700
rect 10832 20640 10896 20644
rect 10912 20700 10976 20704
rect 10912 20644 10916 20700
rect 10916 20644 10972 20700
rect 10972 20644 10976 20700
rect 10912 20640 10976 20644
rect 10992 20700 11056 20704
rect 10992 20644 10996 20700
rect 10996 20644 11052 20700
rect 11052 20644 11056 20700
rect 10992 20640 11056 20644
rect 13752 20700 13816 20704
rect 13752 20644 13756 20700
rect 13756 20644 13812 20700
rect 13812 20644 13816 20700
rect 13752 20640 13816 20644
rect 13832 20700 13896 20704
rect 13832 20644 13836 20700
rect 13836 20644 13892 20700
rect 13892 20644 13896 20700
rect 13832 20640 13896 20644
rect 13912 20700 13976 20704
rect 13912 20644 13916 20700
rect 13916 20644 13972 20700
rect 13972 20644 13976 20700
rect 13912 20640 13976 20644
rect 13992 20700 14056 20704
rect 13992 20644 13996 20700
rect 13996 20644 14052 20700
rect 14052 20644 14056 20700
rect 13992 20640 14056 20644
rect 16752 20700 16816 20704
rect 16752 20644 16756 20700
rect 16756 20644 16812 20700
rect 16812 20644 16816 20700
rect 16752 20640 16816 20644
rect 16832 20700 16896 20704
rect 16832 20644 16836 20700
rect 16836 20644 16892 20700
rect 16892 20644 16896 20700
rect 16832 20640 16896 20644
rect 16912 20700 16976 20704
rect 16912 20644 16916 20700
rect 16916 20644 16972 20700
rect 16972 20644 16976 20700
rect 16912 20640 16976 20644
rect 16992 20700 17056 20704
rect 16992 20644 16996 20700
rect 16996 20644 17052 20700
rect 17052 20644 17056 20700
rect 16992 20640 17056 20644
rect 19752 20700 19816 20704
rect 19752 20644 19756 20700
rect 19756 20644 19812 20700
rect 19812 20644 19816 20700
rect 19752 20640 19816 20644
rect 19832 20700 19896 20704
rect 19832 20644 19836 20700
rect 19836 20644 19892 20700
rect 19892 20644 19896 20700
rect 19832 20640 19896 20644
rect 19912 20700 19976 20704
rect 19912 20644 19916 20700
rect 19916 20644 19972 20700
rect 19972 20644 19976 20700
rect 19912 20640 19976 20644
rect 19992 20700 20056 20704
rect 19992 20644 19996 20700
rect 19996 20644 20052 20700
rect 20052 20644 20056 20700
rect 19992 20640 20056 20644
rect 22752 20700 22816 20704
rect 22752 20644 22756 20700
rect 22756 20644 22812 20700
rect 22812 20644 22816 20700
rect 22752 20640 22816 20644
rect 22832 20700 22896 20704
rect 22832 20644 22836 20700
rect 22836 20644 22892 20700
rect 22892 20644 22896 20700
rect 22832 20640 22896 20644
rect 22912 20700 22976 20704
rect 22912 20644 22916 20700
rect 22916 20644 22972 20700
rect 22972 20644 22976 20700
rect 22912 20640 22976 20644
rect 22992 20700 23056 20704
rect 22992 20644 22996 20700
rect 22996 20644 23052 20700
rect 23052 20644 23056 20700
rect 22992 20640 23056 20644
rect 25752 20700 25816 20704
rect 25752 20644 25756 20700
rect 25756 20644 25812 20700
rect 25812 20644 25816 20700
rect 25752 20640 25816 20644
rect 25832 20700 25896 20704
rect 25832 20644 25836 20700
rect 25836 20644 25892 20700
rect 25892 20644 25896 20700
rect 25832 20640 25896 20644
rect 25912 20700 25976 20704
rect 25912 20644 25916 20700
rect 25916 20644 25972 20700
rect 25972 20644 25976 20700
rect 25912 20640 25976 20644
rect 25992 20700 26056 20704
rect 25992 20644 25996 20700
rect 25996 20644 26052 20700
rect 26052 20644 26056 20700
rect 25992 20640 26056 20644
rect 3252 20156 3316 20160
rect 3252 20100 3256 20156
rect 3256 20100 3312 20156
rect 3312 20100 3316 20156
rect 3252 20096 3316 20100
rect 3332 20156 3396 20160
rect 3332 20100 3336 20156
rect 3336 20100 3392 20156
rect 3392 20100 3396 20156
rect 3332 20096 3396 20100
rect 3412 20156 3476 20160
rect 3412 20100 3416 20156
rect 3416 20100 3472 20156
rect 3472 20100 3476 20156
rect 3412 20096 3476 20100
rect 3492 20156 3556 20160
rect 3492 20100 3496 20156
rect 3496 20100 3552 20156
rect 3552 20100 3556 20156
rect 3492 20096 3556 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 6412 20156 6476 20160
rect 6412 20100 6416 20156
rect 6416 20100 6472 20156
rect 6472 20100 6476 20156
rect 6412 20096 6476 20100
rect 6492 20156 6556 20160
rect 6492 20100 6496 20156
rect 6496 20100 6552 20156
rect 6552 20100 6556 20156
rect 6492 20096 6556 20100
rect 9252 20156 9316 20160
rect 9252 20100 9256 20156
rect 9256 20100 9312 20156
rect 9312 20100 9316 20156
rect 9252 20096 9316 20100
rect 9332 20156 9396 20160
rect 9332 20100 9336 20156
rect 9336 20100 9392 20156
rect 9392 20100 9396 20156
rect 9332 20096 9396 20100
rect 9412 20156 9476 20160
rect 9412 20100 9416 20156
rect 9416 20100 9472 20156
rect 9472 20100 9476 20156
rect 9412 20096 9476 20100
rect 9492 20156 9556 20160
rect 9492 20100 9496 20156
rect 9496 20100 9552 20156
rect 9552 20100 9556 20156
rect 9492 20096 9556 20100
rect 12252 20156 12316 20160
rect 12252 20100 12256 20156
rect 12256 20100 12312 20156
rect 12312 20100 12316 20156
rect 12252 20096 12316 20100
rect 12332 20156 12396 20160
rect 12332 20100 12336 20156
rect 12336 20100 12392 20156
rect 12392 20100 12396 20156
rect 12332 20096 12396 20100
rect 12412 20156 12476 20160
rect 12412 20100 12416 20156
rect 12416 20100 12472 20156
rect 12472 20100 12476 20156
rect 12412 20096 12476 20100
rect 12492 20156 12556 20160
rect 12492 20100 12496 20156
rect 12496 20100 12552 20156
rect 12552 20100 12556 20156
rect 12492 20096 12556 20100
rect 15252 20156 15316 20160
rect 15252 20100 15256 20156
rect 15256 20100 15312 20156
rect 15312 20100 15316 20156
rect 15252 20096 15316 20100
rect 15332 20156 15396 20160
rect 15332 20100 15336 20156
rect 15336 20100 15392 20156
rect 15392 20100 15396 20156
rect 15332 20096 15396 20100
rect 15412 20156 15476 20160
rect 15412 20100 15416 20156
rect 15416 20100 15472 20156
rect 15472 20100 15476 20156
rect 15412 20096 15476 20100
rect 15492 20156 15556 20160
rect 15492 20100 15496 20156
rect 15496 20100 15552 20156
rect 15552 20100 15556 20156
rect 15492 20096 15556 20100
rect 18252 20156 18316 20160
rect 18252 20100 18256 20156
rect 18256 20100 18312 20156
rect 18312 20100 18316 20156
rect 18252 20096 18316 20100
rect 18332 20156 18396 20160
rect 18332 20100 18336 20156
rect 18336 20100 18392 20156
rect 18392 20100 18396 20156
rect 18332 20096 18396 20100
rect 18412 20156 18476 20160
rect 18412 20100 18416 20156
rect 18416 20100 18472 20156
rect 18472 20100 18476 20156
rect 18412 20096 18476 20100
rect 18492 20156 18556 20160
rect 18492 20100 18496 20156
rect 18496 20100 18552 20156
rect 18552 20100 18556 20156
rect 18492 20096 18556 20100
rect 21252 20156 21316 20160
rect 21252 20100 21256 20156
rect 21256 20100 21312 20156
rect 21312 20100 21316 20156
rect 21252 20096 21316 20100
rect 21332 20156 21396 20160
rect 21332 20100 21336 20156
rect 21336 20100 21392 20156
rect 21392 20100 21396 20156
rect 21332 20096 21396 20100
rect 21412 20156 21476 20160
rect 21412 20100 21416 20156
rect 21416 20100 21472 20156
rect 21472 20100 21476 20156
rect 21412 20096 21476 20100
rect 21492 20156 21556 20160
rect 21492 20100 21496 20156
rect 21496 20100 21552 20156
rect 21552 20100 21556 20156
rect 21492 20096 21556 20100
rect 24252 20156 24316 20160
rect 24252 20100 24256 20156
rect 24256 20100 24312 20156
rect 24312 20100 24316 20156
rect 24252 20096 24316 20100
rect 24332 20156 24396 20160
rect 24332 20100 24336 20156
rect 24336 20100 24392 20156
rect 24392 20100 24396 20156
rect 24332 20096 24396 20100
rect 24412 20156 24476 20160
rect 24412 20100 24416 20156
rect 24416 20100 24472 20156
rect 24472 20100 24476 20156
rect 24412 20096 24476 20100
rect 24492 20156 24556 20160
rect 24492 20100 24496 20156
rect 24496 20100 24552 20156
rect 24552 20100 24556 20156
rect 24492 20096 24556 20100
rect 27252 20156 27316 20160
rect 27252 20100 27256 20156
rect 27256 20100 27312 20156
rect 27312 20100 27316 20156
rect 27252 20096 27316 20100
rect 27332 20156 27396 20160
rect 27332 20100 27336 20156
rect 27336 20100 27392 20156
rect 27392 20100 27396 20156
rect 27332 20096 27396 20100
rect 27412 20156 27476 20160
rect 27412 20100 27416 20156
rect 27416 20100 27472 20156
rect 27472 20100 27476 20156
rect 27412 20096 27476 20100
rect 27492 20156 27556 20160
rect 27492 20100 27496 20156
rect 27496 20100 27552 20156
rect 27552 20100 27556 20156
rect 27492 20096 27556 20100
rect 1752 19612 1816 19616
rect 1752 19556 1756 19612
rect 1756 19556 1812 19612
rect 1812 19556 1816 19612
rect 1752 19552 1816 19556
rect 1832 19612 1896 19616
rect 1832 19556 1836 19612
rect 1836 19556 1892 19612
rect 1892 19556 1896 19612
rect 1832 19552 1896 19556
rect 1912 19612 1976 19616
rect 1912 19556 1916 19612
rect 1916 19556 1972 19612
rect 1972 19556 1976 19612
rect 1912 19552 1976 19556
rect 1992 19612 2056 19616
rect 1992 19556 1996 19612
rect 1996 19556 2052 19612
rect 2052 19556 2056 19612
rect 1992 19552 2056 19556
rect 4752 19612 4816 19616
rect 4752 19556 4756 19612
rect 4756 19556 4812 19612
rect 4812 19556 4816 19612
rect 4752 19552 4816 19556
rect 4832 19612 4896 19616
rect 4832 19556 4836 19612
rect 4836 19556 4892 19612
rect 4892 19556 4896 19612
rect 4832 19552 4896 19556
rect 4912 19612 4976 19616
rect 4912 19556 4916 19612
rect 4916 19556 4972 19612
rect 4972 19556 4976 19612
rect 4912 19552 4976 19556
rect 4992 19612 5056 19616
rect 4992 19556 4996 19612
rect 4996 19556 5052 19612
rect 5052 19556 5056 19612
rect 4992 19552 5056 19556
rect 7752 19612 7816 19616
rect 7752 19556 7756 19612
rect 7756 19556 7812 19612
rect 7812 19556 7816 19612
rect 7752 19552 7816 19556
rect 7832 19612 7896 19616
rect 7832 19556 7836 19612
rect 7836 19556 7892 19612
rect 7892 19556 7896 19612
rect 7832 19552 7896 19556
rect 7912 19612 7976 19616
rect 7912 19556 7916 19612
rect 7916 19556 7972 19612
rect 7972 19556 7976 19612
rect 7912 19552 7976 19556
rect 7992 19612 8056 19616
rect 7992 19556 7996 19612
rect 7996 19556 8052 19612
rect 8052 19556 8056 19612
rect 7992 19552 8056 19556
rect 10752 19612 10816 19616
rect 10752 19556 10756 19612
rect 10756 19556 10812 19612
rect 10812 19556 10816 19612
rect 10752 19552 10816 19556
rect 10832 19612 10896 19616
rect 10832 19556 10836 19612
rect 10836 19556 10892 19612
rect 10892 19556 10896 19612
rect 10832 19552 10896 19556
rect 10912 19612 10976 19616
rect 10912 19556 10916 19612
rect 10916 19556 10972 19612
rect 10972 19556 10976 19612
rect 10912 19552 10976 19556
rect 10992 19612 11056 19616
rect 10992 19556 10996 19612
rect 10996 19556 11052 19612
rect 11052 19556 11056 19612
rect 10992 19552 11056 19556
rect 13752 19612 13816 19616
rect 13752 19556 13756 19612
rect 13756 19556 13812 19612
rect 13812 19556 13816 19612
rect 13752 19552 13816 19556
rect 13832 19612 13896 19616
rect 13832 19556 13836 19612
rect 13836 19556 13892 19612
rect 13892 19556 13896 19612
rect 13832 19552 13896 19556
rect 13912 19612 13976 19616
rect 13912 19556 13916 19612
rect 13916 19556 13972 19612
rect 13972 19556 13976 19612
rect 13912 19552 13976 19556
rect 13992 19612 14056 19616
rect 13992 19556 13996 19612
rect 13996 19556 14052 19612
rect 14052 19556 14056 19612
rect 13992 19552 14056 19556
rect 16752 19612 16816 19616
rect 16752 19556 16756 19612
rect 16756 19556 16812 19612
rect 16812 19556 16816 19612
rect 16752 19552 16816 19556
rect 16832 19612 16896 19616
rect 16832 19556 16836 19612
rect 16836 19556 16892 19612
rect 16892 19556 16896 19612
rect 16832 19552 16896 19556
rect 16912 19612 16976 19616
rect 16912 19556 16916 19612
rect 16916 19556 16972 19612
rect 16972 19556 16976 19612
rect 16912 19552 16976 19556
rect 16992 19612 17056 19616
rect 16992 19556 16996 19612
rect 16996 19556 17052 19612
rect 17052 19556 17056 19612
rect 16992 19552 17056 19556
rect 19752 19612 19816 19616
rect 19752 19556 19756 19612
rect 19756 19556 19812 19612
rect 19812 19556 19816 19612
rect 19752 19552 19816 19556
rect 19832 19612 19896 19616
rect 19832 19556 19836 19612
rect 19836 19556 19892 19612
rect 19892 19556 19896 19612
rect 19832 19552 19896 19556
rect 19912 19612 19976 19616
rect 19912 19556 19916 19612
rect 19916 19556 19972 19612
rect 19972 19556 19976 19612
rect 19912 19552 19976 19556
rect 19992 19612 20056 19616
rect 19992 19556 19996 19612
rect 19996 19556 20052 19612
rect 20052 19556 20056 19612
rect 19992 19552 20056 19556
rect 22752 19612 22816 19616
rect 22752 19556 22756 19612
rect 22756 19556 22812 19612
rect 22812 19556 22816 19612
rect 22752 19552 22816 19556
rect 22832 19612 22896 19616
rect 22832 19556 22836 19612
rect 22836 19556 22892 19612
rect 22892 19556 22896 19612
rect 22832 19552 22896 19556
rect 22912 19612 22976 19616
rect 22912 19556 22916 19612
rect 22916 19556 22972 19612
rect 22972 19556 22976 19612
rect 22912 19552 22976 19556
rect 22992 19612 23056 19616
rect 22992 19556 22996 19612
rect 22996 19556 23052 19612
rect 23052 19556 23056 19612
rect 22992 19552 23056 19556
rect 25752 19612 25816 19616
rect 25752 19556 25756 19612
rect 25756 19556 25812 19612
rect 25812 19556 25816 19612
rect 25752 19552 25816 19556
rect 25832 19612 25896 19616
rect 25832 19556 25836 19612
rect 25836 19556 25892 19612
rect 25892 19556 25896 19612
rect 25832 19552 25896 19556
rect 25912 19612 25976 19616
rect 25912 19556 25916 19612
rect 25916 19556 25972 19612
rect 25972 19556 25976 19612
rect 25912 19552 25976 19556
rect 25992 19612 26056 19616
rect 25992 19556 25996 19612
rect 25996 19556 26052 19612
rect 26052 19556 26056 19612
rect 25992 19552 26056 19556
rect 3252 19068 3316 19072
rect 3252 19012 3256 19068
rect 3256 19012 3312 19068
rect 3312 19012 3316 19068
rect 3252 19008 3316 19012
rect 3332 19068 3396 19072
rect 3332 19012 3336 19068
rect 3336 19012 3392 19068
rect 3392 19012 3396 19068
rect 3332 19008 3396 19012
rect 3412 19068 3476 19072
rect 3412 19012 3416 19068
rect 3416 19012 3472 19068
rect 3472 19012 3476 19068
rect 3412 19008 3476 19012
rect 3492 19068 3556 19072
rect 3492 19012 3496 19068
rect 3496 19012 3552 19068
rect 3552 19012 3556 19068
rect 3492 19008 3556 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 6412 19068 6476 19072
rect 6412 19012 6416 19068
rect 6416 19012 6472 19068
rect 6472 19012 6476 19068
rect 6412 19008 6476 19012
rect 6492 19068 6556 19072
rect 6492 19012 6496 19068
rect 6496 19012 6552 19068
rect 6552 19012 6556 19068
rect 6492 19008 6556 19012
rect 9252 19068 9316 19072
rect 9252 19012 9256 19068
rect 9256 19012 9312 19068
rect 9312 19012 9316 19068
rect 9252 19008 9316 19012
rect 9332 19068 9396 19072
rect 9332 19012 9336 19068
rect 9336 19012 9392 19068
rect 9392 19012 9396 19068
rect 9332 19008 9396 19012
rect 9412 19068 9476 19072
rect 9412 19012 9416 19068
rect 9416 19012 9472 19068
rect 9472 19012 9476 19068
rect 9412 19008 9476 19012
rect 9492 19068 9556 19072
rect 9492 19012 9496 19068
rect 9496 19012 9552 19068
rect 9552 19012 9556 19068
rect 9492 19008 9556 19012
rect 12252 19068 12316 19072
rect 12252 19012 12256 19068
rect 12256 19012 12312 19068
rect 12312 19012 12316 19068
rect 12252 19008 12316 19012
rect 12332 19068 12396 19072
rect 12332 19012 12336 19068
rect 12336 19012 12392 19068
rect 12392 19012 12396 19068
rect 12332 19008 12396 19012
rect 12412 19068 12476 19072
rect 12412 19012 12416 19068
rect 12416 19012 12472 19068
rect 12472 19012 12476 19068
rect 12412 19008 12476 19012
rect 12492 19068 12556 19072
rect 12492 19012 12496 19068
rect 12496 19012 12552 19068
rect 12552 19012 12556 19068
rect 12492 19008 12556 19012
rect 15252 19068 15316 19072
rect 15252 19012 15256 19068
rect 15256 19012 15312 19068
rect 15312 19012 15316 19068
rect 15252 19008 15316 19012
rect 15332 19068 15396 19072
rect 15332 19012 15336 19068
rect 15336 19012 15392 19068
rect 15392 19012 15396 19068
rect 15332 19008 15396 19012
rect 15412 19068 15476 19072
rect 15412 19012 15416 19068
rect 15416 19012 15472 19068
rect 15472 19012 15476 19068
rect 15412 19008 15476 19012
rect 15492 19068 15556 19072
rect 15492 19012 15496 19068
rect 15496 19012 15552 19068
rect 15552 19012 15556 19068
rect 15492 19008 15556 19012
rect 18252 19068 18316 19072
rect 18252 19012 18256 19068
rect 18256 19012 18312 19068
rect 18312 19012 18316 19068
rect 18252 19008 18316 19012
rect 18332 19068 18396 19072
rect 18332 19012 18336 19068
rect 18336 19012 18392 19068
rect 18392 19012 18396 19068
rect 18332 19008 18396 19012
rect 18412 19068 18476 19072
rect 18412 19012 18416 19068
rect 18416 19012 18472 19068
rect 18472 19012 18476 19068
rect 18412 19008 18476 19012
rect 18492 19068 18556 19072
rect 18492 19012 18496 19068
rect 18496 19012 18552 19068
rect 18552 19012 18556 19068
rect 18492 19008 18556 19012
rect 21252 19068 21316 19072
rect 21252 19012 21256 19068
rect 21256 19012 21312 19068
rect 21312 19012 21316 19068
rect 21252 19008 21316 19012
rect 21332 19068 21396 19072
rect 21332 19012 21336 19068
rect 21336 19012 21392 19068
rect 21392 19012 21396 19068
rect 21332 19008 21396 19012
rect 21412 19068 21476 19072
rect 21412 19012 21416 19068
rect 21416 19012 21472 19068
rect 21472 19012 21476 19068
rect 21412 19008 21476 19012
rect 21492 19068 21556 19072
rect 21492 19012 21496 19068
rect 21496 19012 21552 19068
rect 21552 19012 21556 19068
rect 21492 19008 21556 19012
rect 24252 19068 24316 19072
rect 24252 19012 24256 19068
rect 24256 19012 24312 19068
rect 24312 19012 24316 19068
rect 24252 19008 24316 19012
rect 24332 19068 24396 19072
rect 24332 19012 24336 19068
rect 24336 19012 24392 19068
rect 24392 19012 24396 19068
rect 24332 19008 24396 19012
rect 24412 19068 24476 19072
rect 24412 19012 24416 19068
rect 24416 19012 24472 19068
rect 24472 19012 24476 19068
rect 24412 19008 24476 19012
rect 24492 19068 24556 19072
rect 24492 19012 24496 19068
rect 24496 19012 24552 19068
rect 24552 19012 24556 19068
rect 24492 19008 24556 19012
rect 27252 19068 27316 19072
rect 27252 19012 27256 19068
rect 27256 19012 27312 19068
rect 27312 19012 27316 19068
rect 27252 19008 27316 19012
rect 27332 19068 27396 19072
rect 27332 19012 27336 19068
rect 27336 19012 27392 19068
rect 27392 19012 27396 19068
rect 27332 19008 27396 19012
rect 27412 19068 27476 19072
rect 27412 19012 27416 19068
rect 27416 19012 27472 19068
rect 27472 19012 27476 19068
rect 27412 19008 27476 19012
rect 27492 19068 27556 19072
rect 27492 19012 27496 19068
rect 27496 19012 27552 19068
rect 27552 19012 27556 19068
rect 27492 19008 27556 19012
rect 1752 18524 1816 18528
rect 1752 18468 1756 18524
rect 1756 18468 1812 18524
rect 1812 18468 1816 18524
rect 1752 18464 1816 18468
rect 1832 18524 1896 18528
rect 1832 18468 1836 18524
rect 1836 18468 1892 18524
rect 1892 18468 1896 18524
rect 1832 18464 1896 18468
rect 1912 18524 1976 18528
rect 1912 18468 1916 18524
rect 1916 18468 1972 18524
rect 1972 18468 1976 18524
rect 1912 18464 1976 18468
rect 1992 18524 2056 18528
rect 1992 18468 1996 18524
rect 1996 18468 2052 18524
rect 2052 18468 2056 18524
rect 1992 18464 2056 18468
rect 4752 18524 4816 18528
rect 4752 18468 4756 18524
rect 4756 18468 4812 18524
rect 4812 18468 4816 18524
rect 4752 18464 4816 18468
rect 4832 18524 4896 18528
rect 4832 18468 4836 18524
rect 4836 18468 4892 18524
rect 4892 18468 4896 18524
rect 4832 18464 4896 18468
rect 4912 18524 4976 18528
rect 4912 18468 4916 18524
rect 4916 18468 4972 18524
rect 4972 18468 4976 18524
rect 4912 18464 4976 18468
rect 4992 18524 5056 18528
rect 4992 18468 4996 18524
rect 4996 18468 5052 18524
rect 5052 18468 5056 18524
rect 4992 18464 5056 18468
rect 7752 18524 7816 18528
rect 7752 18468 7756 18524
rect 7756 18468 7812 18524
rect 7812 18468 7816 18524
rect 7752 18464 7816 18468
rect 7832 18524 7896 18528
rect 7832 18468 7836 18524
rect 7836 18468 7892 18524
rect 7892 18468 7896 18524
rect 7832 18464 7896 18468
rect 7912 18524 7976 18528
rect 7912 18468 7916 18524
rect 7916 18468 7972 18524
rect 7972 18468 7976 18524
rect 7912 18464 7976 18468
rect 7992 18524 8056 18528
rect 7992 18468 7996 18524
rect 7996 18468 8052 18524
rect 8052 18468 8056 18524
rect 7992 18464 8056 18468
rect 10752 18524 10816 18528
rect 10752 18468 10756 18524
rect 10756 18468 10812 18524
rect 10812 18468 10816 18524
rect 10752 18464 10816 18468
rect 10832 18524 10896 18528
rect 10832 18468 10836 18524
rect 10836 18468 10892 18524
rect 10892 18468 10896 18524
rect 10832 18464 10896 18468
rect 10912 18524 10976 18528
rect 10912 18468 10916 18524
rect 10916 18468 10972 18524
rect 10972 18468 10976 18524
rect 10912 18464 10976 18468
rect 10992 18524 11056 18528
rect 10992 18468 10996 18524
rect 10996 18468 11052 18524
rect 11052 18468 11056 18524
rect 10992 18464 11056 18468
rect 13752 18524 13816 18528
rect 13752 18468 13756 18524
rect 13756 18468 13812 18524
rect 13812 18468 13816 18524
rect 13752 18464 13816 18468
rect 13832 18524 13896 18528
rect 13832 18468 13836 18524
rect 13836 18468 13892 18524
rect 13892 18468 13896 18524
rect 13832 18464 13896 18468
rect 13912 18524 13976 18528
rect 13912 18468 13916 18524
rect 13916 18468 13972 18524
rect 13972 18468 13976 18524
rect 13912 18464 13976 18468
rect 13992 18524 14056 18528
rect 13992 18468 13996 18524
rect 13996 18468 14052 18524
rect 14052 18468 14056 18524
rect 13992 18464 14056 18468
rect 16752 18524 16816 18528
rect 16752 18468 16756 18524
rect 16756 18468 16812 18524
rect 16812 18468 16816 18524
rect 16752 18464 16816 18468
rect 16832 18524 16896 18528
rect 16832 18468 16836 18524
rect 16836 18468 16892 18524
rect 16892 18468 16896 18524
rect 16832 18464 16896 18468
rect 16912 18524 16976 18528
rect 16912 18468 16916 18524
rect 16916 18468 16972 18524
rect 16972 18468 16976 18524
rect 16912 18464 16976 18468
rect 16992 18524 17056 18528
rect 16992 18468 16996 18524
rect 16996 18468 17052 18524
rect 17052 18468 17056 18524
rect 16992 18464 17056 18468
rect 19752 18524 19816 18528
rect 19752 18468 19756 18524
rect 19756 18468 19812 18524
rect 19812 18468 19816 18524
rect 19752 18464 19816 18468
rect 19832 18524 19896 18528
rect 19832 18468 19836 18524
rect 19836 18468 19892 18524
rect 19892 18468 19896 18524
rect 19832 18464 19896 18468
rect 19912 18524 19976 18528
rect 19912 18468 19916 18524
rect 19916 18468 19972 18524
rect 19972 18468 19976 18524
rect 19912 18464 19976 18468
rect 19992 18524 20056 18528
rect 19992 18468 19996 18524
rect 19996 18468 20052 18524
rect 20052 18468 20056 18524
rect 19992 18464 20056 18468
rect 22752 18524 22816 18528
rect 22752 18468 22756 18524
rect 22756 18468 22812 18524
rect 22812 18468 22816 18524
rect 22752 18464 22816 18468
rect 22832 18524 22896 18528
rect 22832 18468 22836 18524
rect 22836 18468 22892 18524
rect 22892 18468 22896 18524
rect 22832 18464 22896 18468
rect 22912 18524 22976 18528
rect 22912 18468 22916 18524
rect 22916 18468 22972 18524
rect 22972 18468 22976 18524
rect 22912 18464 22976 18468
rect 22992 18524 23056 18528
rect 22992 18468 22996 18524
rect 22996 18468 23052 18524
rect 23052 18468 23056 18524
rect 22992 18464 23056 18468
rect 25752 18524 25816 18528
rect 25752 18468 25756 18524
rect 25756 18468 25812 18524
rect 25812 18468 25816 18524
rect 25752 18464 25816 18468
rect 25832 18524 25896 18528
rect 25832 18468 25836 18524
rect 25836 18468 25892 18524
rect 25892 18468 25896 18524
rect 25832 18464 25896 18468
rect 25912 18524 25976 18528
rect 25912 18468 25916 18524
rect 25916 18468 25972 18524
rect 25972 18468 25976 18524
rect 25912 18464 25976 18468
rect 25992 18524 26056 18528
rect 25992 18468 25996 18524
rect 25996 18468 26052 18524
rect 26052 18468 26056 18524
rect 25992 18464 26056 18468
rect 3252 17980 3316 17984
rect 3252 17924 3256 17980
rect 3256 17924 3312 17980
rect 3312 17924 3316 17980
rect 3252 17920 3316 17924
rect 3332 17980 3396 17984
rect 3332 17924 3336 17980
rect 3336 17924 3392 17980
rect 3392 17924 3396 17980
rect 3332 17920 3396 17924
rect 3412 17980 3476 17984
rect 3412 17924 3416 17980
rect 3416 17924 3472 17980
rect 3472 17924 3476 17980
rect 3412 17920 3476 17924
rect 3492 17980 3556 17984
rect 3492 17924 3496 17980
rect 3496 17924 3552 17980
rect 3552 17924 3556 17980
rect 3492 17920 3556 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 6412 17980 6476 17984
rect 6412 17924 6416 17980
rect 6416 17924 6472 17980
rect 6472 17924 6476 17980
rect 6412 17920 6476 17924
rect 6492 17980 6556 17984
rect 6492 17924 6496 17980
rect 6496 17924 6552 17980
rect 6552 17924 6556 17980
rect 6492 17920 6556 17924
rect 9252 17980 9316 17984
rect 9252 17924 9256 17980
rect 9256 17924 9312 17980
rect 9312 17924 9316 17980
rect 9252 17920 9316 17924
rect 9332 17980 9396 17984
rect 9332 17924 9336 17980
rect 9336 17924 9392 17980
rect 9392 17924 9396 17980
rect 9332 17920 9396 17924
rect 9412 17980 9476 17984
rect 9412 17924 9416 17980
rect 9416 17924 9472 17980
rect 9472 17924 9476 17980
rect 9412 17920 9476 17924
rect 9492 17980 9556 17984
rect 9492 17924 9496 17980
rect 9496 17924 9552 17980
rect 9552 17924 9556 17980
rect 9492 17920 9556 17924
rect 12252 17980 12316 17984
rect 12252 17924 12256 17980
rect 12256 17924 12312 17980
rect 12312 17924 12316 17980
rect 12252 17920 12316 17924
rect 12332 17980 12396 17984
rect 12332 17924 12336 17980
rect 12336 17924 12392 17980
rect 12392 17924 12396 17980
rect 12332 17920 12396 17924
rect 12412 17980 12476 17984
rect 12412 17924 12416 17980
rect 12416 17924 12472 17980
rect 12472 17924 12476 17980
rect 12412 17920 12476 17924
rect 12492 17980 12556 17984
rect 12492 17924 12496 17980
rect 12496 17924 12552 17980
rect 12552 17924 12556 17980
rect 12492 17920 12556 17924
rect 15252 17980 15316 17984
rect 15252 17924 15256 17980
rect 15256 17924 15312 17980
rect 15312 17924 15316 17980
rect 15252 17920 15316 17924
rect 15332 17980 15396 17984
rect 15332 17924 15336 17980
rect 15336 17924 15392 17980
rect 15392 17924 15396 17980
rect 15332 17920 15396 17924
rect 15412 17980 15476 17984
rect 15412 17924 15416 17980
rect 15416 17924 15472 17980
rect 15472 17924 15476 17980
rect 15412 17920 15476 17924
rect 15492 17980 15556 17984
rect 15492 17924 15496 17980
rect 15496 17924 15552 17980
rect 15552 17924 15556 17980
rect 15492 17920 15556 17924
rect 18252 17980 18316 17984
rect 18252 17924 18256 17980
rect 18256 17924 18312 17980
rect 18312 17924 18316 17980
rect 18252 17920 18316 17924
rect 18332 17980 18396 17984
rect 18332 17924 18336 17980
rect 18336 17924 18392 17980
rect 18392 17924 18396 17980
rect 18332 17920 18396 17924
rect 18412 17980 18476 17984
rect 18412 17924 18416 17980
rect 18416 17924 18472 17980
rect 18472 17924 18476 17980
rect 18412 17920 18476 17924
rect 18492 17980 18556 17984
rect 18492 17924 18496 17980
rect 18496 17924 18552 17980
rect 18552 17924 18556 17980
rect 18492 17920 18556 17924
rect 21252 17980 21316 17984
rect 21252 17924 21256 17980
rect 21256 17924 21312 17980
rect 21312 17924 21316 17980
rect 21252 17920 21316 17924
rect 21332 17980 21396 17984
rect 21332 17924 21336 17980
rect 21336 17924 21392 17980
rect 21392 17924 21396 17980
rect 21332 17920 21396 17924
rect 21412 17980 21476 17984
rect 21412 17924 21416 17980
rect 21416 17924 21472 17980
rect 21472 17924 21476 17980
rect 21412 17920 21476 17924
rect 21492 17980 21556 17984
rect 21492 17924 21496 17980
rect 21496 17924 21552 17980
rect 21552 17924 21556 17980
rect 21492 17920 21556 17924
rect 24252 17980 24316 17984
rect 24252 17924 24256 17980
rect 24256 17924 24312 17980
rect 24312 17924 24316 17980
rect 24252 17920 24316 17924
rect 24332 17980 24396 17984
rect 24332 17924 24336 17980
rect 24336 17924 24392 17980
rect 24392 17924 24396 17980
rect 24332 17920 24396 17924
rect 24412 17980 24476 17984
rect 24412 17924 24416 17980
rect 24416 17924 24472 17980
rect 24472 17924 24476 17980
rect 24412 17920 24476 17924
rect 24492 17980 24556 17984
rect 24492 17924 24496 17980
rect 24496 17924 24552 17980
rect 24552 17924 24556 17980
rect 24492 17920 24556 17924
rect 27252 17980 27316 17984
rect 27252 17924 27256 17980
rect 27256 17924 27312 17980
rect 27312 17924 27316 17980
rect 27252 17920 27316 17924
rect 27332 17980 27396 17984
rect 27332 17924 27336 17980
rect 27336 17924 27392 17980
rect 27392 17924 27396 17980
rect 27332 17920 27396 17924
rect 27412 17980 27476 17984
rect 27412 17924 27416 17980
rect 27416 17924 27472 17980
rect 27472 17924 27476 17980
rect 27412 17920 27476 17924
rect 27492 17980 27556 17984
rect 27492 17924 27496 17980
rect 27496 17924 27552 17980
rect 27552 17924 27556 17980
rect 27492 17920 27556 17924
rect 1752 17436 1816 17440
rect 1752 17380 1756 17436
rect 1756 17380 1812 17436
rect 1812 17380 1816 17436
rect 1752 17376 1816 17380
rect 1832 17436 1896 17440
rect 1832 17380 1836 17436
rect 1836 17380 1892 17436
rect 1892 17380 1896 17436
rect 1832 17376 1896 17380
rect 1912 17436 1976 17440
rect 1912 17380 1916 17436
rect 1916 17380 1972 17436
rect 1972 17380 1976 17436
rect 1912 17376 1976 17380
rect 1992 17436 2056 17440
rect 1992 17380 1996 17436
rect 1996 17380 2052 17436
rect 2052 17380 2056 17436
rect 1992 17376 2056 17380
rect 4752 17436 4816 17440
rect 4752 17380 4756 17436
rect 4756 17380 4812 17436
rect 4812 17380 4816 17436
rect 4752 17376 4816 17380
rect 4832 17436 4896 17440
rect 4832 17380 4836 17436
rect 4836 17380 4892 17436
rect 4892 17380 4896 17436
rect 4832 17376 4896 17380
rect 4912 17436 4976 17440
rect 4912 17380 4916 17436
rect 4916 17380 4972 17436
rect 4972 17380 4976 17436
rect 4912 17376 4976 17380
rect 4992 17436 5056 17440
rect 4992 17380 4996 17436
rect 4996 17380 5052 17436
rect 5052 17380 5056 17436
rect 4992 17376 5056 17380
rect 7752 17436 7816 17440
rect 7752 17380 7756 17436
rect 7756 17380 7812 17436
rect 7812 17380 7816 17436
rect 7752 17376 7816 17380
rect 7832 17436 7896 17440
rect 7832 17380 7836 17436
rect 7836 17380 7892 17436
rect 7892 17380 7896 17436
rect 7832 17376 7896 17380
rect 7912 17436 7976 17440
rect 7912 17380 7916 17436
rect 7916 17380 7972 17436
rect 7972 17380 7976 17436
rect 7912 17376 7976 17380
rect 7992 17436 8056 17440
rect 7992 17380 7996 17436
rect 7996 17380 8052 17436
rect 8052 17380 8056 17436
rect 7992 17376 8056 17380
rect 10752 17436 10816 17440
rect 10752 17380 10756 17436
rect 10756 17380 10812 17436
rect 10812 17380 10816 17436
rect 10752 17376 10816 17380
rect 10832 17436 10896 17440
rect 10832 17380 10836 17436
rect 10836 17380 10892 17436
rect 10892 17380 10896 17436
rect 10832 17376 10896 17380
rect 10912 17436 10976 17440
rect 10912 17380 10916 17436
rect 10916 17380 10972 17436
rect 10972 17380 10976 17436
rect 10912 17376 10976 17380
rect 10992 17436 11056 17440
rect 10992 17380 10996 17436
rect 10996 17380 11052 17436
rect 11052 17380 11056 17436
rect 10992 17376 11056 17380
rect 13752 17436 13816 17440
rect 13752 17380 13756 17436
rect 13756 17380 13812 17436
rect 13812 17380 13816 17436
rect 13752 17376 13816 17380
rect 13832 17436 13896 17440
rect 13832 17380 13836 17436
rect 13836 17380 13892 17436
rect 13892 17380 13896 17436
rect 13832 17376 13896 17380
rect 13912 17436 13976 17440
rect 13912 17380 13916 17436
rect 13916 17380 13972 17436
rect 13972 17380 13976 17436
rect 13912 17376 13976 17380
rect 13992 17436 14056 17440
rect 13992 17380 13996 17436
rect 13996 17380 14052 17436
rect 14052 17380 14056 17436
rect 13992 17376 14056 17380
rect 16752 17436 16816 17440
rect 16752 17380 16756 17436
rect 16756 17380 16812 17436
rect 16812 17380 16816 17436
rect 16752 17376 16816 17380
rect 16832 17436 16896 17440
rect 16832 17380 16836 17436
rect 16836 17380 16892 17436
rect 16892 17380 16896 17436
rect 16832 17376 16896 17380
rect 16912 17436 16976 17440
rect 16912 17380 16916 17436
rect 16916 17380 16972 17436
rect 16972 17380 16976 17436
rect 16912 17376 16976 17380
rect 16992 17436 17056 17440
rect 16992 17380 16996 17436
rect 16996 17380 17052 17436
rect 17052 17380 17056 17436
rect 16992 17376 17056 17380
rect 19752 17436 19816 17440
rect 19752 17380 19756 17436
rect 19756 17380 19812 17436
rect 19812 17380 19816 17436
rect 19752 17376 19816 17380
rect 19832 17436 19896 17440
rect 19832 17380 19836 17436
rect 19836 17380 19892 17436
rect 19892 17380 19896 17436
rect 19832 17376 19896 17380
rect 19912 17436 19976 17440
rect 19912 17380 19916 17436
rect 19916 17380 19972 17436
rect 19972 17380 19976 17436
rect 19912 17376 19976 17380
rect 19992 17436 20056 17440
rect 19992 17380 19996 17436
rect 19996 17380 20052 17436
rect 20052 17380 20056 17436
rect 19992 17376 20056 17380
rect 22752 17436 22816 17440
rect 22752 17380 22756 17436
rect 22756 17380 22812 17436
rect 22812 17380 22816 17436
rect 22752 17376 22816 17380
rect 22832 17436 22896 17440
rect 22832 17380 22836 17436
rect 22836 17380 22892 17436
rect 22892 17380 22896 17436
rect 22832 17376 22896 17380
rect 22912 17436 22976 17440
rect 22912 17380 22916 17436
rect 22916 17380 22972 17436
rect 22972 17380 22976 17436
rect 22912 17376 22976 17380
rect 22992 17436 23056 17440
rect 22992 17380 22996 17436
rect 22996 17380 23052 17436
rect 23052 17380 23056 17436
rect 22992 17376 23056 17380
rect 25752 17436 25816 17440
rect 25752 17380 25756 17436
rect 25756 17380 25812 17436
rect 25812 17380 25816 17436
rect 25752 17376 25816 17380
rect 25832 17436 25896 17440
rect 25832 17380 25836 17436
rect 25836 17380 25892 17436
rect 25892 17380 25896 17436
rect 25832 17376 25896 17380
rect 25912 17436 25976 17440
rect 25912 17380 25916 17436
rect 25916 17380 25972 17436
rect 25972 17380 25976 17436
rect 25912 17376 25976 17380
rect 25992 17436 26056 17440
rect 25992 17380 25996 17436
rect 25996 17380 26052 17436
rect 26052 17380 26056 17436
rect 25992 17376 26056 17380
rect 3252 16892 3316 16896
rect 3252 16836 3256 16892
rect 3256 16836 3312 16892
rect 3312 16836 3316 16892
rect 3252 16832 3316 16836
rect 3332 16892 3396 16896
rect 3332 16836 3336 16892
rect 3336 16836 3392 16892
rect 3392 16836 3396 16892
rect 3332 16832 3396 16836
rect 3412 16892 3476 16896
rect 3412 16836 3416 16892
rect 3416 16836 3472 16892
rect 3472 16836 3476 16892
rect 3412 16832 3476 16836
rect 3492 16892 3556 16896
rect 3492 16836 3496 16892
rect 3496 16836 3552 16892
rect 3552 16836 3556 16892
rect 3492 16832 3556 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 6412 16892 6476 16896
rect 6412 16836 6416 16892
rect 6416 16836 6472 16892
rect 6472 16836 6476 16892
rect 6412 16832 6476 16836
rect 6492 16892 6556 16896
rect 6492 16836 6496 16892
rect 6496 16836 6552 16892
rect 6552 16836 6556 16892
rect 6492 16832 6556 16836
rect 9252 16892 9316 16896
rect 9252 16836 9256 16892
rect 9256 16836 9312 16892
rect 9312 16836 9316 16892
rect 9252 16832 9316 16836
rect 9332 16892 9396 16896
rect 9332 16836 9336 16892
rect 9336 16836 9392 16892
rect 9392 16836 9396 16892
rect 9332 16832 9396 16836
rect 9412 16892 9476 16896
rect 9412 16836 9416 16892
rect 9416 16836 9472 16892
rect 9472 16836 9476 16892
rect 9412 16832 9476 16836
rect 9492 16892 9556 16896
rect 9492 16836 9496 16892
rect 9496 16836 9552 16892
rect 9552 16836 9556 16892
rect 9492 16832 9556 16836
rect 12252 16892 12316 16896
rect 12252 16836 12256 16892
rect 12256 16836 12312 16892
rect 12312 16836 12316 16892
rect 12252 16832 12316 16836
rect 12332 16892 12396 16896
rect 12332 16836 12336 16892
rect 12336 16836 12392 16892
rect 12392 16836 12396 16892
rect 12332 16832 12396 16836
rect 12412 16892 12476 16896
rect 12412 16836 12416 16892
rect 12416 16836 12472 16892
rect 12472 16836 12476 16892
rect 12412 16832 12476 16836
rect 12492 16892 12556 16896
rect 12492 16836 12496 16892
rect 12496 16836 12552 16892
rect 12552 16836 12556 16892
rect 12492 16832 12556 16836
rect 15252 16892 15316 16896
rect 15252 16836 15256 16892
rect 15256 16836 15312 16892
rect 15312 16836 15316 16892
rect 15252 16832 15316 16836
rect 15332 16892 15396 16896
rect 15332 16836 15336 16892
rect 15336 16836 15392 16892
rect 15392 16836 15396 16892
rect 15332 16832 15396 16836
rect 15412 16892 15476 16896
rect 15412 16836 15416 16892
rect 15416 16836 15472 16892
rect 15472 16836 15476 16892
rect 15412 16832 15476 16836
rect 15492 16892 15556 16896
rect 15492 16836 15496 16892
rect 15496 16836 15552 16892
rect 15552 16836 15556 16892
rect 15492 16832 15556 16836
rect 18252 16892 18316 16896
rect 18252 16836 18256 16892
rect 18256 16836 18312 16892
rect 18312 16836 18316 16892
rect 18252 16832 18316 16836
rect 18332 16892 18396 16896
rect 18332 16836 18336 16892
rect 18336 16836 18392 16892
rect 18392 16836 18396 16892
rect 18332 16832 18396 16836
rect 18412 16892 18476 16896
rect 18412 16836 18416 16892
rect 18416 16836 18472 16892
rect 18472 16836 18476 16892
rect 18412 16832 18476 16836
rect 18492 16892 18556 16896
rect 18492 16836 18496 16892
rect 18496 16836 18552 16892
rect 18552 16836 18556 16892
rect 18492 16832 18556 16836
rect 21252 16892 21316 16896
rect 21252 16836 21256 16892
rect 21256 16836 21312 16892
rect 21312 16836 21316 16892
rect 21252 16832 21316 16836
rect 21332 16892 21396 16896
rect 21332 16836 21336 16892
rect 21336 16836 21392 16892
rect 21392 16836 21396 16892
rect 21332 16832 21396 16836
rect 21412 16892 21476 16896
rect 21412 16836 21416 16892
rect 21416 16836 21472 16892
rect 21472 16836 21476 16892
rect 21412 16832 21476 16836
rect 21492 16892 21556 16896
rect 21492 16836 21496 16892
rect 21496 16836 21552 16892
rect 21552 16836 21556 16892
rect 21492 16832 21556 16836
rect 24252 16892 24316 16896
rect 24252 16836 24256 16892
rect 24256 16836 24312 16892
rect 24312 16836 24316 16892
rect 24252 16832 24316 16836
rect 24332 16892 24396 16896
rect 24332 16836 24336 16892
rect 24336 16836 24392 16892
rect 24392 16836 24396 16892
rect 24332 16832 24396 16836
rect 24412 16892 24476 16896
rect 24412 16836 24416 16892
rect 24416 16836 24472 16892
rect 24472 16836 24476 16892
rect 24412 16832 24476 16836
rect 24492 16892 24556 16896
rect 24492 16836 24496 16892
rect 24496 16836 24552 16892
rect 24552 16836 24556 16892
rect 24492 16832 24556 16836
rect 27252 16892 27316 16896
rect 27252 16836 27256 16892
rect 27256 16836 27312 16892
rect 27312 16836 27316 16892
rect 27252 16832 27316 16836
rect 27332 16892 27396 16896
rect 27332 16836 27336 16892
rect 27336 16836 27392 16892
rect 27392 16836 27396 16892
rect 27332 16832 27396 16836
rect 27412 16892 27476 16896
rect 27412 16836 27416 16892
rect 27416 16836 27472 16892
rect 27472 16836 27476 16892
rect 27412 16832 27476 16836
rect 27492 16892 27556 16896
rect 27492 16836 27496 16892
rect 27496 16836 27552 16892
rect 27552 16836 27556 16892
rect 27492 16832 27556 16836
rect 1752 16348 1816 16352
rect 1752 16292 1756 16348
rect 1756 16292 1812 16348
rect 1812 16292 1816 16348
rect 1752 16288 1816 16292
rect 1832 16348 1896 16352
rect 1832 16292 1836 16348
rect 1836 16292 1892 16348
rect 1892 16292 1896 16348
rect 1832 16288 1896 16292
rect 1912 16348 1976 16352
rect 1912 16292 1916 16348
rect 1916 16292 1972 16348
rect 1972 16292 1976 16348
rect 1912 16288 1976 16292
rect 1992 16348 2056 16352
rect 1992 16292 1996 16348
rect 1996 16292 2052 16348
rect 2052 16292 2056 16348
rect 1992 16288 2056 16292
rect 4752 16348 4816 16352
rect 4752 16292 4756 16348
rect 4756 16292 4812 16348
rect 4812 16292 4816 16348
rect 4752 16288 4816 16292
rect 4832 16348 4896 16352
rect 4832 16292 4836 16348
rect 4836 16292 4892 16348
rect 4892 16292 4896 16348
rect 4832 16288 4896 16292
rect 4912 16348 4976 16352
rect 4912 16292 4916 16348
rect 4916 16292 4972 16348
rect 4972 16292 4976 16348
rect 4912 16288 4976 16292
rect 4992 16348 5056 16352
rect 4992 16292 4996 16348
rect 4996 16292 5052 16348
rect 5052 16292 5056 16348
rect 4992 16288 5056 16292
rect 7752 16348 7816 16352
rect 7752 16292 7756 16348
rect 7756 16292 7812 16348
rect 7812 16292 7816 16348
rect 7752 16288 7816 16292
rect 7832 16348 7896 16352
rect 7832 16292 7836 16348
rect 7836 16292 7892 16348
rect 7892 16292 7896 16348
rect 7832 16288 7896 16292
rect 7912 16348 7976 16352
rect 7912 16292 7916 16348
rect 7916 16292 7972 16348
rect 7972 16292 7976 16348
rect 7912 16288 7976 16292
rect 7992 16348 8056 16352
rect 7992 16292 7996 16348
rect 7996 16292 8052 16348
rect 8052 16292 8056 16348
rect 7992 16288 8056 16292
rect 10752 16348 10816 16352
rect 10752 16292 10756 16348
rect 10756 16292 10812 16348
rect 10812 16292 10816 16348
rect 10752 16288 10816 16292
rect 10832 16348 10896 16352
rect 10832 16292 10836 16348
rect 10836 16292 10892 16348
rect 10892 16292 10896 16348
rect 10832 16288 10896 16292
rect 10912 16348 10976 16352
rect 10912 16292 10916 16348
rect 10916 16292 10972 16348
rect 10972 16292 10976 16348
rect 10912 16288 10976 16292
rect 10992 16348 11056 16352
rect 10992 16292 10996 16348
rect 10996 16292 11052 16348
rect 11052 16292 11056 16348
rect 10992 16288 11056 16292
rect 13752 16348 13816 16352
rect 13752 16292 13756 16348
rect 13756 16292 13812 16348
rect 13812 16292 13816 16348
rect 13752 16288 13816 16292
rect 13832 16348 13896 16352
rect 13832 16292 13836 16348
rect 13836 16292 13892 16348
rect 13892 16292 13896 16348
rect 13832 16288 13896 16292
rect 13912 16348 13976 16352
rect 13912 16292 13916 16348
rect 13916 16292 13972 16348
rect 13972 16292 13976 16348
rect 13912 16288 13976 16292
rect 13992 16348 14056 16352
rect 13992 16292 13996 16348
rect 13996 16292 14052 16348
rect 14052 16292 14056 16348
rect 13992 16288 14056 16292
rect 16752 16348 16816 16352
rect 16752 16292 16756 16348
rect 16756 16292 16812 16348
rect 16812 16292 16816 16348
rect 16752 16288 16816 16292
rect 16832 16348 16896 16352
rect 16832 16292 16836 16348
rect 16836 16292 16892 16348
rect 16892 16292 16896 16348
rect 16832 16288 16896 16292
rect 16912 16348 16976 16352
rect 16912 16292 16916 16348
rect 16916 16292 16972 16348
rect 16972 16292 16976 16348
rect 16912 16288 16976 16292
rect 16992 16348 17056 16352
rect 16992 16292 16996 16348
rect 16996 16292 17052 16348
rect 17052 16292 17056 16348
rect 16992 16288 17056 16292
rect 19752 16348 19816 16352
rect 19752 16292 19756 16348
rect 19756 16292 19812 16348
rect 19812 16292 19816 16348
rect 19752 16288 19816 16292
rect 19832 16348 19896 16352
rect 19832 16292 19836 16348
rect 19836 16292 19892 16348
rect 19892 16292 19896 16348
rect 19832 16288 19896 16292
rect 19912 16348 19976 16352
rect 19912 16292 19916 16348
rect 19916 16292 19972 16348
rect 19972 16292 19976 16348
rect 19912 16288 19976 16292
rect 19992 16348 20056 16352
rect 19992 16292 19996 16348
rect 19996 16292 20052 16348
rect 20052 16292 20056 16348
rect 19992 16288 20056 16292
rect 22752 16348 22816 16352
rect 22752 16292 22756 16348
rect 22756 16292 22812 16348
rect 22812 16292 22816 16348
rect 22752 16288 22816 16292
rect 22832 16348 22896 16352
rect 22832 16292 22836 16348
rect 22836 16292 22892 16348
rect 22892 16292 22896 16348
rect 22832 16288 22896 16292
rect 22912 16348 22976 16352
rect 22912 16292 22916 16348
rect 22916 16292 22972 16348
rect 22972 16292 22976 16348
rect 22912 16288 22976 16292
rect 22992 16348 23056 16352
rect 22992 16292 22996 16348
rect 22996 16292 23052 16348
rect 23052 16292 23056 16348
rect 22992 16288 23056 16292
rect 25752 16348 25816 16352
rect 25752 16292 25756 16348
rect 25756 16292 25812 16348
rect 25812 16292 25816 16348
rect 25752 16288 25816 16292
rect 25832 16348 25896 16352
rect 25832 16292 25836 16348
rect 25836 16292 25892 16348
rect 25892 16292 25896 16348
rect 25832 16288 25896 16292
rect 25912 16348 25976 16352
rect 25912 16292 25916 16348
rect 25916 16292 25972 16348
rect 25972 16292 25976 16348
rect 25912 16288 25976 16292
rect 25992 16348 26056 16352
rect 25992 16292 25996 16348
rect 25996 16292 26052 16348
rect 26052 16292 26056 16348
rect 25992 16288 26056 16292
rect 3252 15804 3316 15808
rect 3252 15748 3256 15804
rect 3256 15748 3312 15804
rect 3312 15748 3316 15804
rect 3252 15744 3316 15748
rect 3332 15804 3396 15808
rect 3332 15748 3336 15804
rect 3336 15748 3392 15804
rect 3392 15748 3396 15804
rect 3332 15744 3396 15748
rect 3412 15804 3476 15808
rect 3412 15748 3416 15804
rect 3416 15748 3472 15804
rect 3472 15748 3476 15804
rect 3412 15744 3476 15748
rect 3492 15804 3556 15808
rect 3492 15748 3496 15804
rect 3496 15748 3552 15804
rect 3552 15748 3556 15804
rect 3492 15744 3556 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 6412 15804 6476 15808
rect 6412 15748 6416 15804
rect 6416 15748 6472 15804
rect 6472 15748 6476 15804
rect 6412 15744 6476 15748
rect 6492 15804 6556 15808
rect 6492 15748 6496 15804
rect 6496 15748 6552 15804
rect 6552 15748 6556 15804
rect 6492 15744 6556 15748
rect 9252 15804 9316 15808
rect 9252 15748 9256 15804
rect 9256 15748 9312 15804
rect 9312 15748 9316 15804
rect 9252 15744 9316 15748
rect 9332 15804 9396 15808
rect 9332 15748 9336 15804
rect 9336 15748 9392 15804
rect 9392 15748 9396 15804
rect 9332 15744 9396 15748
rect 9412 15804 9476 15808
rect 9412 15748 9416 15804
rect 9416 15748 9472 15804
rect 9472 15748 9476 15804
rect 9412 15744 9476 15748
rect 9492 15804 9556 15808
rect 9492 15748 9496 15804
rect 9496 15748 9552 15804
rect 9552 15748 9556 15804
rect 9492 15744 9556 15748
rect 12252 15804 12316 15808
rect 12252 15748 12256 15804
rect 12256 15748 12312 15804
rect 12312 15748 12316 15804
rect 12252 15744 12316 15748
rect 12332 15804 12396 15808
rect 12332 15748 12336 15804
rect 12336 15748 12392 15804
rect 12392 15748 12396 15804
rect 12332 15744 12396 15748
rect 12412 15804 12476 15808
rect 12412 15748 12416 15804
rect 12416 15748 12472 15804
rect 12472 15748 12476 15804
rect 12412 15744 12476 15748
rect 12492 15804 12556 15808
rect 12492 15748 12496 15804
rect 12496 15748 12552 15804
rect 12552 15748 12556 15804
rect 12492 15744 12556 15748
rect 15252 15804 15316 15808
rect 15252 15748 15256 15804
rect 15256 15748 15312 15804
rect 15312 15748 15316 15804
rect 15252 15744 15316 15748
rect 15332 15804 15396 15808
rect 15332 15748 15336 15804
rect 15336 15748 15392 15804
rect 15392 15748 15396 15804
rect 15332 15744 15396 15748
rect 15412 15804 15476 15808
rect 15412 15748 15416 15804
rect 15416 15748 15472 15804
rect 15472 15748 15476 15804
rect 15412 15744 15476 15748
rect 15492 15804 15556 15808
rect 15492 15748 15496 15804
rect 15496 15748 15552 15804
rect 15552 15748 15556 15804
rect 15492 15744 15556 15748
rect 18252 15804 18316 15808
rect 18252 15748 18256 15804
rect 18256 15748 18312 15804
rect 18312 15748 18316 15804
rect 18252 15744 18316 15748
rect 18332 15804 18396 15808
rect 18332 15748 18336 15804
rect 18336 15748 18392 15804
rect 18392 15748 18396 15804
rect 18332 15744 18396 15748
rect 18412 15804 18476 15808
rect 18412 15748 18416 15804
rect 18416 15748 18472 15804
rect 18472 15748 18476 15804
rect 18412 15744 18476 15748
rect 18492 15804 18556 15808
rect 18492 15748 18496 15804
rect 18496 15748 18552 15804
rect 18552 15748 18556 15804
rect 18492 15744 18556 15748
rect 21252 15804 21316 15808
rect 21252 15748 21256 15804
rect 21256 15748 21312 15804
rect 21312 15748 21316 15804
rect 21252 15744 21316 15748
rect 21332 15804 21396 15808
rect 21332 15748 21336 15804
rect 21336 15748 21392 15804
rect 21392 15748 21396 15804
rect 21332 15744 21396 15748
rect 21412 15804 21476 15808
rect 21412 15748 21416 15804
rect 21416 15748 21472 15804
rect 21472 15748 21476 15804
rect 21412 15744 21476 15748
rect 21492 15804 21556 15808
rect 21492 15748 21496 15804
rect 21496 15748 21552 15804
rect 21552 15748 21556 15804
rect 21492 15744 21556 15748
rect 24252 15804 24316 15808
rect 24252 15748 24256 15804
rect 24256 15748 24312 15804
rect 24312 15748 24316 15804
rect 24252 15744 24316 15748
rect 24332 15804 24396 15808
rect 24332 15748 24336 15804
rect 24336 15748 24392 15804
rect 24392 15748 24396 15804
rect 24332 15744 24396 15748
rect 24412 15804 24476 15808
rect 24412 15748 24416 15804
rect 24416 15748 24472 15804
rect 24472 15748 24476 15804
rect 24412 15744 24476 15748
rect 24492 15804 24556 15808
rect 24492 15748 24496 15804
rect 24496 15748 24552 15804
rect 24552 15748 24556 15804
rect 24492 15744 24556 15748
rect 27252 15804 27316 15808
rect 27252 15748 27256 15804
rect 27256 15748 27312 15804
rect 27312 15748 27316 15804
rect 27252 15744 27316 15748
rect 27332 15804 27396 15808
rect 27332 15748 27336 15804
rect 27336 15748 27392 15804
rect 27392 15748 27396 15804
rect 27332 15744 27396 15748
rect 27412 15804 27476 15808
rect 27412 15748 27416 15804
rect 27416 15748 27472 15804
rect 27472 15748 27476 15804
rect 27412 15744 27476 15748
rect 27492 15804 27556 15808
rect 27492 15748 27496 15804
rect 27496 15748 27552 15804
rect 27552 15748 27556 15804
rect 27492 15744 27556 15748
rect 1752 15260 1816 15264
rect 1752 15204 1756 15260
rect 1756 15204 1812 15260
rect 1812 15204 1816 15260
rect 1752 15200 1816 15204
rect 1832 15260 1896 15264
rect 1832 15204 1836 15260
rect 1836 15204 1892 15260
rect 1892 15204 1896 15260
rect 1832 15200 1896 15204
rect 1912 15260 1976 15264
rect 1912 15204 1916 15260
rect 1916 15204 1972 15260
rect 1972 15204 1976 15260
rect 1912 15200 1976 15204
rect 1992 15260 2056 15264
rect 1992 15204 1996 15260
rect 1996 15204 2052 15260
rect 2052 15204 2056 15260
rect 1992 15200 2056 15204
rect 4752 15260 4816 15264
rect 4752 15204 4756 15260
rect 4756 15204 4812 15260
rect 4812 15204 4816 15260
rect 4752 15200 4816 15204
rect 4832 15260 4896 15264
rect 4832 15204 4836 15260
rect 4836 15204 4892 15260
rect 4892 15204 4896 15260
rect 4832 15200 4896 15204
rect 4912 15260 4976 15264
rect 4912 15204 4916 15260
rect 4916 15204 4972 15260
rect 4972 15204 4976 15260
rect 4912 15200 4976 15204
rect 4992 15260 5056 15264
rect 4992 15204 4996 15260
rect 4996 15204 5052 15260
rect 5052 15204 5056 15260
rect 4992 15200 5056 15204
rect 7752 15260 7816 15264
rect 7752 15204 7756 15260
rect 7756 15204 7812 15260
rect 7812 15204 7816 15260
rect 7752 15200 7816 15204
rect 7832 15260 7896 15264
rect 7832 15204 7836 15260
rect 7836 15204 7892 15260
rect 7892 15204 7896 15260
rect 7832 15200 7896 15204
rect 7912 15260 7976 15264
rect 7912 15204 7916 15260
rect 7916 15204 7972 15260
rect 7972 15204 7976 15260
rect 7912 15200 7976 15204
rect 7992 15260 8056 15264
rect 7992 15204 7996 15260
rect 7996 15204 8052 15260
rect 8052 15204 8056 15260
rect 7992 15200 8056 15204
rect 10752 15260 10816 15264
rect 10752 15204 10756 15260
rect 10756 15204 10812 15260
rect 10812 15204 10816 15260
rect 10752 15200 10816 15204
rect 10832 15260 10896 15264
rect 10832 15204 10836 15260
rect 10836 15204 10892 15260
rect 10892 15204 10896 15260
rect 10832 15200 10896 15204
rect 10912 15260 10976 15264
rect 10912 15204 10916 15260
rect 10916 15204 10972 15260
rect 10972 15204 10976 15260
rect 10912 15200 10976 15204
rect 10992 15260 11056 15264
rect 10992 15204 10996 15260
rect 10996 15204 11052 15260
rect 11052 15204 11056 15260
rect 10992 15200 11056 15204
rect 13752 15260 13816 15264
rect 13752 15204 13756 15260
rect 13756 15204 13812 15260
rect 13812 15204 13816 15260
rect 13752 15200 13816 15204
rect 13832 15260 13896 15264
rect 13832 15204 13836 15260
rect 13836 15204 13892 15260
rect 13892 15204 13896 15260
rect 13832 15200 13896 15204
rect 13912 15260 13976 15264
rect 13912 15204 13916 15260
rect 13916 15204 13972 15260
rect 13972 15204 13976 15260
rect 13912 15200 13976 15204
rect 13992 15260 14056 15264
rect 13992 15204 13996 15260
rect 13996 15204 14052 15260
rect 14052 15204 14056 15260
rect 13992 15200 14056 15204
rect 16752 15260 16816 15264
rect 16752 15204 16756 15260
rect 16756 15204 16812 15260
rect 16812 15204 16816 15260
rect 16752 15200 16816 15204
rect 16832 15260 16896 15264
rect 16832 15204 16836 15260
rect 16836 15204 16892 15260
rect 16892 15204 16896 15260
rect 16832 15200 16896 15204
rect 16912 15260 16976 15264
rect 16912 15204 16916 15260
rect 16916 15204 16972 15260
rect 16972 15204 16976 15260
rect 16912 15200 16976 15204
rect 16992 15260 17056 15264
rect 16992 15204 16996 15260
rect 16996 15204 17052 15260
rect 17052 15204 17056 15260
rect 16992 15200 17056 15204
rect 19752 15260 19816 15264
rect 19752 15204 19756 15260
rect 19756 15204 19812 15260
rect 19812 15204 19816 15260
rect 19752 15200 19816 15204
rect 19832 15260 19896 15264
rect 19832 15204 19836 15260
rect 19836 15204 19892 15260
rect 19892 15204 19896 15260
rect 19832 15200 19896 15204
rect 19912 15260 19976 15264
rect 19912 15204 19916 15260
rect 19916 15204 19972 15260
rect 19972 15204 19976 15260
rect 19912 15200 19976 15204
rect 19992 15260 20056 15264
rect 19992 15204 19996 15260
rect 19996 15204 20052 15260
rect 20052 15204 20056 15260
rect 19992 15200 20056 15204
rect 22752 15260 22816 15264
rect 22752 15204 22756 15260
rect 22756 15204 22812 15260
rect 22812 15204 22816 15260
rect 22752 15200 22816 15204
rect 22832 15260 22896 15264
rect 22832 15204 22836 15260
rect 22836 15204 22892 15260
rect 22892 15204 22896 15260
rect 22832 15200 22896 15204
rect 22912 15260 22976 15264
rect 22912 15204 22916 15260
rect 22916 15204 22972 15260
rect 22972 15204 22976 15260
rect 22912 15200 22976 15204
rect 22992 15260 23056 15264
rect 22992 15204 22996 15260
rect 22996 15204 23052 15260
rect 23052 15204 23056 15260
rect 22992 15200 23056 15204
rect 25752 15260 25816 15264
rect 25752 15204 25756 15260
rect 25756 15204 25812 15260
rect 25812 15204 25816 15260
rect 25752 15200 25816 15204
rect 25832 15260 25896 15264
rect 25832 15204 25836 15260
rect 25836 15204 25892 15260
rect 25892 15204 25896 15260
rect 25832 15200 25896 15204
rect 25912 15260 25976 15264
rect 25912 15204 25916 15260
rect 25916 15204 25972 15260
rect 25972 15204 25976 15260
rect 25912 15200 25976 15204
rect 25992 15260 26056 15264
rect 25992 15204 25996 15260
rect 25996 15204 26052 15260
rect 26052 15204 26056 15260
rect 25992 15200 26056 15204
rect 3252 14716 3316 14720
rect 3252 14660 3256 14716
rect 3256 14660 3312 14716
rect 3312 14660 3316 14716
rect 3252 14656 3316 14660
rect 3332 14716 3396 14720
rect 3332 14660 3336 14716
rect 3336 14660 3392 14716
rect 3392 14660 3396 14716
rect 3332 14656 3396 14660
rect 3412 14716 3476 14720
rect 3412 14660 3416 14716
rect 3416 14660 3472 14716
rect 3472 14660 3476 14716
rect 3412 14656 3476 14660
rect 3492 14716 3556 14720
rect 3492 14660 3496 14716
rect 3496 14660 3552 14716
rect 3552 14660 3556 14716
rect 3492 14656 3556 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 6412 14716 6476 14720
rect 6412 14660 6416 14716
rect 6416 14660 6472 14716
rect 6472 14660 6476 14716
rect 6412 14656 6476 14660
rect 6492 14716 6556 14720
rect 6492 14660 6496 14716
rect 6496 14660 6552 14716
rect 6552 14660 6556 14716
rect 6492 14656 6556 14660
rect 9252 14716 9316 14720
rect 9252 14660 9256 14716
rect 9256 14660 9312 14716
rect 9312 14660 9316 14716
rect 9252 14656 9316 14660
rect 9332 14716 9396 14720
rect 9332 14660 9336 14716
rect 9336 14660 9392 14716
rect 9392 14660 9396 14716
rect 9332 14656 9396 14660
rect 9412 14716 9476 14720
rect 9412 14660 9416 14716
rect 9416 14660 9472 14716
rect 9472 14660 9476 14716
rect 9412 14656 9476 14660
rect 9492 14716 9556 14720
rect 9492 14660 9496 14716
rect 9496 14660 9552 14716
rect 9552 14660 9556 14716
rect 9492 14656 9556 14660
rect 12252 14716 12316 14720
rect 12252 14660 12256 14716
rect 12256 14660 12312 14716
rect 12312 14660 12316 14716
rect 12252 14656 12316 14660
rect 12332 14716 12396 14720
rect 12332 14660 12336 14716
rect 12336 14660 12392 14716
rect 12392 14660 12396 14716
rect 12332 14656 12396 14660
rect 12412 14716 12476 14720
rect 12412 14660 12416 14716
rect 12416 14660 12472 14716
rect 12472 14660 12476 14716
rect 12412 14656 12476 14660
rect 12492 14716 12556 14720
rect 12492 14660 12496 14716
rect 12496 14660 12552 14716
rect 12552 14660 12556 14716
rect 12492 14656 12556 14660
rect 15252 14716 15316 14720
rect 15252 14660 15256 14716
rect 15256 14660 15312 14716
rect 15312 14660 15316 14716
rect 15252 14656 15316 14660
rect 15332 14716 15396 14720
rect 15332 14660 15336 14716
rect 15336 14660 15392 14716
rect 15392 14660 15396 14716
rect 15332 14656 15396 14660
rect 15412 14716 15476 14720
rect 15412 14660 15416 14716
rect 15416 14660 15472 14716
rect 15472 14660 15476 14716
rect 15412 14656 15476 14660
rect 15492 14716 15556 14720
rect 15492 14660 15496 14716
rect 15496 14660 15552 14716
rect 15552 14660 15556 14716
rect 15492 14656 15556 14660
rect 18252 14716 18316 14720
rect 18252 14660 18256 14716
rect 18256 14660 18312 14716
rect 18312 14660 18316 14716
rect 18252 14656 18316 14660
rect 18332 14716 18396 14720
rect 18332 14660 18336 14716
rect 18336 14660 18392 14716
rect 18392 14660 18396 14716
rect 18332 14656 18396 14660
rect 18412 14716 18476 14720
rect 18412 14660 18416 14716
rect 18416 14660 18472 14716
rect 18472 14660 18476 14716
rect 18412 14656 18476 14660
rect 18492 14716 18556 14720
rect 18492 14660 18496 14716
rect 18496 14660 18552 14716
rect 18552 14660 18556 14716
rect 18492 14656 18556 14660
rect 21252 14716 21316 14720
rect 21252 14660 21256 14716
rect 21256 14660 21312 14716
rect 21312 14660 21316 14716
rect 21252 14656 21316 14660
rect 21332 14716 21396 14720
rect 21332 14660 21336 14716
rect 21336 14660 21392 14716
rect 21392 14660 21396 14716
rect 21332 14656 21396 14660
rect 21412 14716 21476 14720
rect 21412 14660 21416 14716
rect 21416 14660 21472 14716
rect 21472 14660 21476 14716
rect 21412 14656 21476 14660
rect 21492 14716 21556 14720
rect 21492 14660 21496 14716
rect 21496 14660 21552 14716
rect 21552 14660 21556 14716
rect 21492 14656 21556 14660
rect 24252 14716 24316 14720
rect 24252 14660 24256 14716
rect 24256 14660 24312 14716
rect 24312 14660 24316 14716
rect 24252 14656 24316 14660
rect 24332 14716 24396 14720
rect 24332 14660 24336 14716
rect 24336 14660 24392 14716
rect 24392 14660 24396 14716
rect 24332 14656 24396 14660
rect 24412 14716 24476 14720
rect 24412 14660 24416 14716
rect 24416 14660 24472 14716
rect 24472 14660 24476 14716
rect 24412 14656 24476 14660
rect 24492 14716 24556 14720
rect 24492 14660 24496 14716
rect 24496 14660 24552 14716
rect 24552 14660 24556 14716
rect 24492 14656 24556 14660
rect 27252 14716 27316 14720
rect 27252 14660 27256 14716
rect 27256 14660 27312 14716
rect 27312 14660 27316 14716
rect 27252 14656 27316 14660
rect 27332 14716 27396 14720
rect 27332 14660 27336 14716
rect 27336 14660 27392 14716
rect 27392 14660 27396 14716
rect 27332 14656 27396 14660
rect 27412 14716 27476 14720
rect 27412 14660 27416 14716
rect 27416 14660 27472 14716
rect 27472 14660 27476 14716
rect 27412 14656 27476 14660
rect 27492 14716 27556 14720
rect 27492 14660 27496 14716
rect 27496 14660 27552 14716
rect 27552 14660 27556 14716
rect 27492 14656 27556 14660
rect 1752 14172 1816 14176
rect 1752 14116 1756 14172
rect 1756 14116 1812 14172
rect 1812 14116 1816 14172
rect 1752 14112 1816 14116
rect 1832 14172 1896 14176
rect 1832 14116 1836 14172
rect 1836 14116 1892 14172
rect 1892 14116 1896 14172
rect 1832 14112 1896 14116
rect 1912 14172 1976 14176
rect 1912 14116 1916 14172
rect 1916 14116 1972 14172
rect 1972 14116 1976 14172
rect 1912 14112 1976 14116
rect 1992 14172 2056 14176
rect 1992 14116 1996 14172
rect 1996 14116 2052 14172
rect 2052 14116 2056 14172
rect 1992 14112 2056 14116
rect 4752 14172 4816 14176
rect 4752 14116 4756 14172
rect 4756 14116 4812 14172
rect 4812 14116 4816 14172
rect 4752 14112 4816 14116
rect 4832 14172 4896 14176
rect 4832 14116 4836 14172
rect 4836 14116 4892 14172
rect 4892 14116 4896 14172
rect 4832 14112 4896 14116
rect 4912 14172 4976 14176
rect 4912 14116 4916 14172
rect 4916 14116 4972 14172
rect 4972 14116 4976 14172
rect 4912 14112 4976 14116
rect 4992 14172 5056 14176
rect 4992 14116 4996 14172
rect 4996 14116 5052 14172
rect 5052 14116 5056 14172
rect 4992 14112 5056 14116
rect 7752 14172 7816 14176
rect 7752 14116 7756 14172
rect 7756 14116 7812 14172
rect 7812 14116 7816 14172
rect 7752 14112 7816 14116
rect 7832 14172 7896 14176
rect 7832 14116 7836 14172
rect 7836 14116 7892 14172
rect 7892 14116 7896 14172
rect 7832 14112 7896 14116
rect 7912 14172 7976 14176
rect 7912 14116 7916 14172
rect 7916 14116 7972 14172
rect 7972 14116 7976 14172
rect 7912 14112 7976 14116
rect 7992 14172 8056 14176
rect 7992 14116 7996 14172
rect 7996 14116 8052 14172
rect 8052 14116 8056 14172
rect 7992 14112 8056 14116
rect 10752 14172 10816 14176
rect 10752 14116 10756 14172
rect 10756 14116 10812 14172
rect 10812 14116 10816 14172
rect 10752 14112 10816 14116
rect 10832 14172 10896 14176
rect 10832 14116 10836 14172
rect 10836 14116 10892 14172
rect 10892 14116 10896 14172
rect 10832 14112 10896 14116
rect 10912 14172 10976 14176
rect 10912 14116 10916 14172
rect 10916 14116 10972 14172
rect 10972 14116 10976 14172
rect 10912 14112 10976 14116
rect 10992 14172 11056 14176
rect 10992 14116 10996 14172
rect 10996 14116 11052 14172
rect 11052 14116 11056 14172
rect 10992 14112 11056 14116
rect 13752 14172 13816 14176
rect 13752 14116 13756 14172
rect 13756 14116 13812 14172
rect 13812 14116 13816 14172
rect 13752 14112 13816 14116
rect 13832 14172 13896 14176
rect 13832 14116 13836 14172
rect 13836 14116 13892 14172
rect 13892 14116 13896 14172
rect 13832 14112 13896 14116
rect 13912 14172 13976 14176
rect 13912 14116 13916 14172
rect 13916 14116 13972 14172
rect 13972 14116 13976 14172
rect 13912 14112 13976 14116
rect 13992 14172 14056 14176
rect 13992 14116 13996 14172
rect 13996 14116 14052 14172
rect 14052 14116 14056 14172
rect 13992 14112 14056 14116
rect 16752 14172 16816 14176
rect 16752 14116 16756 14172
rect 16756 14116 16812 14172
rect 16812 14116 16816 14172
rect 16752 14112 16816 14116
rect 16832 14172 16896 14176
rect 16832 14116 16836 14172
rect 16836 14116 16892 14172
rect 16892 14116 16896 14172
rect 16832 14112 16896 14116
rect 16912 14172 16976 14176
rect 16912 14116 16916 14172
rect 16916 14116 16972 14172
rect 16972 14116 16976 14172
rect 16912 14112 16976 14116
rect 16992 14172 17056 14176
rect 16992 14116 16996 14172
rect 16996 14116 17052 14172
rect 17052 14116 17056 14172
rect 16992 14112 17056 14116
rect 19752 14172 19816 14176
rect 19752 14116 19756 14172
rect 19756 14116 19812 14172
rect 19812 14116 19816 14172
rect 19752 14112 19816 14116
rect 19832 14172 19896 14176
rect 19832 14116 19836 14172
rect 19836 14116 19892 14172
rect 19892 14116 19896 14172
rect 19832 14112 19896 14116
rect 19912 14172 19976 14176
rect 19912 14116 19916 14172
rect 19916 14116 19972 14172
rect 19972 14116 19976 14172
rect 19912 14112 19976 14116
rect 19992 14172 20056 14176
rect 19992 14116 19996 14172
rect 19996 14116 20052 14172
rect 20052 14116 20056 14172
rect 19992 14112 20056 14116
rect 22752 14172 22816 14176
rect 22752 14116 22756 14172
rect 22756 14116 22812 14172
rect 22812 14116 22816 14172
rect 22752 14112 22816 14116
rect 22832 14172 22896 14176
rect 22832 14116 22836 14172
rect 22836 14116 22892 14172
rect 22892 14116 22896 14172
rect 22832 14112 22896 14116
rect 22912 14172 22976 14176
rect 22912 14116 22916 14172
rect 22916 14116 22972 14172
rect 22972 14116 22976 14172
rect 22912 14112 22976 14116
rect 22992 14172 23056 14176
rect 22992 14116 22996 14172
rect 22996 14116 23052 14172
rect 23052 14116 23056 14172
rect 22992 14112 23056 14116
rect 25752 14172 25816 14176
rect 25752 14116 25756 14172
rect 25756 14116 25812 14172
rect 25812 14116 25816 14172
rect 25752 14112 25816 14116
rect 25832 14172 25896 14176
rect 25832 14116 25836 14172
rect 25836 14116 25892 14172
rect 25892 14116 25896 14172
rect 25832 14112 25896 14116
rect 25912 14172 25976 14176
rect 25912 14116 25916 14172
rect 25916 14116 25972 14172
rect 25972 14116 25976 14172
rect 25912 14112 25976 14116
rect 25992 14172 26056 14176
rect 25992 14116 25996 14172
rect 25996 14116 26052 14172
rect 26052 14116 26056 14172
rect 25992 14112 26056 14116
rect 3252 13628 3316 13632
rect 3252 13572 3256 13628
rect 3256 13572 3312 13628
rect 3312 13572 3316 13628
rect 3252 13568 3316 13572
rect 3332 13628 3396 13632
rect 3332 13572 3336 13628
rect 3336 13572 3392 13628
rect 3392 13572 3396 13628
rect 3332 13568 3396 13572
rect 3412 13628 3476 13632
rect 3412 13572 3416 13628
rect 3416 13572 3472 13628
rect 3472 13572 3476 13628
rect 3412 13568 3476 13572
rect 3492 13628 3556 13632
rect 3492 13572 3496 13628
rect 3496 13572 3552 13628
rect 3552 13572 3556 13628
rect 3492 13568 3556 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 6412 13628 6476 13632
rect 6412 13572 6416 13628
rect 6416 13572 6472 13628
rect 6472 13572 6476 13628
rect 6412 13568 6476 13572
rect 6492 13628 6556 13632
rect 6492 13572 6496 13628
rect 6496 13572 6552 13628
rect 6552 13572 6556 13628
rect 6492 13568 6556 13572
rect 9252 13628 9316 13632
rect 9252 13572 9256 13628
rect 9256 13572 9312 13628
rect 9312 13572 9316 13628
rect 9252 13568 9316 13572
rect 9332 13628 9396 13632
rect 9332 13572 9336 13628
rect 9336 13572 9392 13628
rect 9392 13572 9396 13628
rect 9332 13568 9396 13572
rect 9412 13628 9476 13632
rect 9412 13572 9416 13628
rect 9416 13572 9472 13628
rect 9472 13572 9476 13628
rect 9412 13568 9476 13572
rect 9492 13628 9556 13632
rect 9492 13572 9496 13628
rect 9496 13572 9552 13628
rect 9552 13572 9556 13628
rect 9492 13568 9556 13572
rect 12252 13628 12316 13632
rect 12252 13572 12256 13628
rect 12256 13572 12312 13628
rect 12312 13572 12316 13628
rect 12252 13568 12316 13572
rect 12332 13628 12396 13632
rect 12332 13572 12336 13628
rect 12336 13572 12392 13628
rect 12392 13572 12396 13628
rect 12332 13568 12396 13572
rect 12412 13628 12476 13632
rect 12412 13572 12416 13628
rect 12416 13572 12472 13628
rect 12472 13572 12476 13628
rect 12412 13568 12476 13572
rect 12492 13628 12556 13632
rect 12492 13572 12496 13628
rect 12496 13572 12552 13628
rect 12552 13572 12556 13628
rect 12492 13568 12556 13572
rect 15252 13628 15316 13632
rect 15252 13572 15256 13628
rect 15256 13572 15312 13628
rect 15312 13572 15316 13628
rect 15252 13568 15316 13572
rect 15332 13628 15396 13632
rect 15332 13572 15336 13628
rect 15336 13572 15392 13628
rect 15392 13572 15396 13628
rect 15332 13568 15396 13572
rect 15412 13628 15476 13632
rect 15412 13572 15416 13628
rect 15416 13572 15472 13628
rect 15472 13572 15476 13628
rect 15412 13568 15476 13572
rect 15492 13628 15556 13632
rect 15492 13572 15496 13628
rect 15496 13572 15552 13628
rect 15552 13572 15556 13628
rect 15492 13568 15556 13572
rect 18252 13628 18316 13632
rect 18252 13572 18256 13628
rect 18256 13572 18312 13628
rect 18312 13572 18316 13628
rect 18252 13568 18316 13572
rect 18332 13628 18396 13632
rect 18332 13572 18336 13628
rect 18336 13572 18392 13628
rect 18392 13572 18396 13628
rect 18332 13568 18396 13572
rect 18412 13628 18476 13632
rect 18412 13572 18416 13628
rect 18416 13572 18472 13628
rect 18472 13572 18476 13628
rect 18412 13568 18476 13572
rect 18492 13628 18556 13632
rect 18492 13572 18496 13628
rect 18496 13572 18552 13628
rect 18552 13572 18556 13628
rect 18492 13568 18556 13572
rect 21252 13628 21316 13632
rect 21252 13572 21256 13628
rect 21256 13572 21312 13628
rect 21312 13572 21316 13628
rect 21252 13568 21316 13572
rect 21332 13628 21396 13632
rect 21332 13572 21336 13628
rect 21336 13572 21392 13628
rect 21392 13572 21396 13628
rect 21332 13568 21396 13572
rect 21412 13628 21476 13632
rect 21412 13572 21416 13628
rect 21416 13572 21472 13628
rect 21472 13572 21476 13628
rect 21412 13568 21476 13572
rect 21492 13628 21556 13632
rect 21492 13572 21496 13628
rect 21496 13572 21552 13628
rect 21552 13572 21556 13628
rect 21492 13568 21556 13572
rect 24252 13628 24316 13632
rect 24252 13572 24256 13628
rect 24256 13572 24312 13628
rect 24312 13572 24316 13628
rect 24252 13568 24316 13572
rect 24332 13628 24396 13632
rect 24332 13572 24336 13628
rect 24336 13572 24392 13628
rect 24392 13572 24396 13628
rect 24332 13568 24396 13572
rect 24412 13628 24476 13632
rect 24412 13572 24416 13628
rect 24416 13572 24472 13628
rect 24472 13572 24476 13628
rect 24412 13568 24476 13572
rect 24492 13628 24556 13632
rect 24492 13572 24496 13628
rect 24496 13572 24552 13628
rect 24552 13572 24556 13628
rect 24492 13568 24556 13572
rect 27252 13628 27316 13632
rect 27252 13572 27256 13628
rect 27256 13572 27312 13628
rect 27312 13572 27316 13628
rect 27252 13568 27316 13572
rect 27332 13628 27396 13632
rect 27332 13572 27336 13628
rect 27336 13572 27392 13628
rect 27392 13572 27396 13628
rect 27332 13568 27396 13572
rect 27412 13628 27476 13632
rect 27412 13572 27416 13628
rect 27416 13572 27472 13628
rect 27472 13572 27476 13628
rect 27412 13568 27476 13572
rect 27492 13628 27556 13632
rect 27492 13572 27496 13628
rect 27496 13572 27552 13628
rect 27552 13572 27556 13628
rect 27492 13568 27556 13572
rect 1752 13084 1816 13088
rect 1752 13028 1756 13084
rect 1756 13028 1812 13084
rect 1812 13028 1816 13084
rect 1752 13024 1816 13028
rect 1832 13084 1896 13088
rect 1832 13028 1836 13084
rect 1836 13028 1892 13084
rect 1892 13028 1896 13084
rect 1832 13024 1896 13028
rect 1912 13084 1976 13088
rect 1912 13028 1916 13084
rect 1916 13028 1972 13084
rect 1972 13028 1976 13084
rect 1912 13024 1976 13028
rect 1992 13084 2056 13088
rect 1992 13028 1996 13084
rect 1996 13028 2052 13084
rect 2052 13028 2056 13084
rect 1992 13024 2056 13028
rect 4752 13084 4816 13088
rect 4752 13028 4756 13084
rect 4756 13028 4812 13084
rect 4812 13028 4816 13084
rect 4752 13024 4816 13028
rect 4832 13084 4896 13088
rect 4832 13028 4836 13084
rect 4836 13028 4892 13084
rect 4892 13028 4896 13084
rect 4832 13024 4896 13028
rect 4912 13084 4976 13088
rect 4912 13028 4916 13084
rect 4916 13028 4972 13084
rect 4972 13028 4976 13084
rect 4912 13024 4976 13028
rect 4992 13084 5056 13088
rect 4992 13028 4996 13084
rect 4996 13028 5052 13084
rect 5052 13028 5056 13084
rect 4992 13024 5056 13028
rect 7752 13084 7816 13088
rect 7752 13028 7756 13084
rect 7756 13028 7812 13084
rect 7812 13028 7816 13084
rect 7752 13024 7816 13028
rect 7832 13084 7896 13088
rect 7832 13028 7836 13084
rect 7836 13028 7892 13084
rect 7892 13028 7896 13084
rect 7832 13024 7896 13028
rect 7912 13084 7976 13088
rect 7912 13028 7916 13084
rect 7916 13028 7972 13084
rect 7972 13028 7976 13084
rect 7912 13024 7976 13028
rect 7992 13084 8056 13088
rect 7992 13028 7996 13084
rect 7996 13028 8052 13084
rect 8052 13028 8056 13084
rect 7992 13024 8056 13028
rect 10752 13084 10816 13088
rect 10752 13028 10756 13084
rect 10756 13028 10812 13084
rect 10812 13028 10816 13084
rect 10752 13024 10816 13028
rect 10832 13084 10896 13088
rect 10832 13028 10836 13084
rect 10836 13028 10892 13084
rect 10892 13028 10896 13084
rect 10832 13024 10896 13028
rect 10912 13084 10976 13088
rect 10912 13028 10916 13084
rect 10916 13028 10972 13084
rect 10972 13028 10976 13084
rect 10912 13024 10976 13028
rect 10992 13084 11056 13088
rect 10992 13028 10996 13084
rect 10996 13028 11052 13084
rect 11052 13028 11056 13084
rect 10992 13024 11056 13028
rect 13752 13084 13816 13088
rect 13752 13028 13756 13084
rect 13756 13028 13812 13084
rect 13812 13028 13816 13084
rect 13752 13024 13816 13028
rect 13832 13084 13896 13088
rect 13832 13028 13836 13084
rect 13836 13028 13892 13084
rect 13892 13028 13896 13084
rect 13832 13024 13896 13028
rect 13912 13084 13976 13088
rect 13912 13028 13916 13084
rect 13916 13028 13972 13084
rect 13972 13028 13976 13084
rect 13912 13024 13976 13028
rect 13992 13084 14056 13088
rect 13992 13028 13996 13084
rect 13996 13028 14052 13084
rect 14052 13028 14056 13084
rect 13992 13024 14056 13028
rect 16752 13084 16816 13088
rect 16752 13028 16756 13084
rect 16756 13028 16812 13084
rect 16812 13028 16816 13084
rect 16752 13024 16816 13028
rect 16832 13084 16896 13088
rect 16832 13028 16836 13084
rect 16836 13028 16892 13084
rect 16892 13028 16896 13084
rect 16832 13024 16896 13028
rect 16912 13084 16976 13088
rect 16912 13028 16916 13084
rect 16916 13028 16972 13084
rect 16972 13028 16976 13084
rect 16912 13024 16976 13028
rect 16992 13084 17056 13088
rect 16992 13028 16996 13084
rect 16996 13028 17052 13084
rect 17052 13028 17056 13084
rect 16992 13024 17056 13028
rect 19752 13084 19816 13088
rect 19752 13028 19756 13084
rect 19756 13028 19812 13084
rect 19812 13028 19816 13084
rect 19752 13024 19816 13028
rect 19832 13084 19896 13088
rect 19832 13028 19836 13084
rect 19836 13028 19892 13084
rect 19892 13028 19896 13084
rect 19832 13024 19896 13028
rect 19912 13084 19976 13088
rect 19912 13028 19916 13084
rect 19916 13028 19972 13084
rect 19972 13028 19976 13084
rect 19912 13024 19976 13028
rect 19992 13084 20056 13088
rect 19992 13028 19996 13084
rect 19996 13028 20052 13084
rect 20052 13028 20056 13084
rect 19992 13024 20056 13028
rect 22752 13084 22816 13088
rect 22752 13028 22756 13084
rect 22756 13028 22812 13084
rect 22812 13028 22816 13084
rect 22752 13024 22816 13028
rect 22832 13084 22896 13088
rect 22832 13028 22836 13084
rect 22836 13028 22892 13084
rect 22892 13028 22896 13084
rect 22832 13024 22896 13028
rect 22912 13084 22976 13088
rect 22912 13028 22916 13084
rect 22916 13028 22972 13084
rect 22972 13028 22976 13084
rect 22912 13024 22976 13028
rect 22992 13084 23056 13088
rect 22992 13028 22996 13084
rect 22996 13028 23052 13084
rect 23052 13028 23056 13084
rect 22992 13024 23056 13028
rect 25752 13084 25816 13088
rect 25752 13028 25756 13084
rect 25756 13028 25812 13084
rect 25812 13028 25816 13084
rect 25752 13024 25816 13028
rect 25832 13084 25896 13088
rect 25832 13028 25836 13084
rect 25836 13028 25892 13084
rect 25892 13028 25896 13084
rect 25832 13024 25896 13028
rect 25912 13084 25976 13088
rect 25912 13028 25916 13084
rect 25916 13028 25972 13084
rect 25972 13028 25976 13084
rect 25912 13024 25976 13028
rect 25992 13084 26056 13088
rect 25992 13028 25996 13084
rect 25996 13028 26052 13084
rect 26052 13028 26056 13084
rect 25992 13024 26056 13028
rect 3252 12540 3316 12544
rect 3252 12484 3256 12540
rect 3256 12484 3312 12540
rect 3312 12484 3316 12540
rect 3252 12480 3316 12484
rect 3332 12540 3396 12544
rect 3332 12484 3336 12540
rect 3336 12484 3392 12540
rect 3392 12484 3396 12540
rect 3332 12480 3396 12484
rect 3412 12540 3476 12544
rect 3412 12484 3416 12540
rect 3416 12484 3472 12540
rect 3472 12484 3476 12540
rect 3412 12480 3476 12484
rect 3492 12540 3556 12544
rect 3492 12484 3496 12540
rect 3496 12484 3552 12540
rect 3552 12484 3556 12540
rect 3492 12480 3556 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 6412 12540 6476 12544
rect 6412 12484 6416 12540
rect 6416 12484 6472 12540
rect 6472 12484 6476 12540
rect 6412 12480 6476 12484
rect 6492 12540 6556 12544
rect 6492 12484 6496 12540
rect 6496 12484 6552 12540
rect 6552 12484 6556 12540
rect 6492 12480 6556 12484
rect 9252 12540 9316 12544
rect 9252 12484 9256 12540
rect 9256 12484 9312 12540
rect 9312 12484 9316 12540
rect 9252 12480 9316 12484
rect 9332 12540 9396 12544
rect 9332 12484 9336 12540
rect 9336 12484 9392 12540
rect 9392 12484 9396 12540
rect 9332 12480 9396 12484
rect 9412 12540 9476 12544
rect 9412 12484 9416 12540
rect 9416 12484 9472 12540
rect 9472 12484 9476 12540
rect 9412 12480 9476 12484
rect 9492 12540 9556 12544
rect 9492 12484 9496 12540
rect 9496 12484 9552 12540
rect 9552 12484 9556 12540
rect 9492 12480 9556 12484
rect 12252 12540 12316 12544
rect 12252 12484 12256 12540
rect 12256 12484 12312 12540
rect 12312 12484 12316 12540
rect 12252 12480 12316 12484
rect 12332 12540 12396 12544
rect 12332 12484 12336 12540
rect 12336 12484 12392 12540
rect 12392 12484 12396 12540
rect 12332 12480 12396 12484
rect 12412 12540 12476 12544
rect 12412 12484 12416 12540
rect 12416 12484 12472 12540
rect 12472 12484 12476 12540
rect 12412 12480 12476 12484
rect 12492 12540 12556 12544
rect 12492 12484 12496 12540
rect 12496 12484 12552 12540
rect 12552 12484 12556 12540
rect 12492 12480 12556 12484
rect 15252 12540 15316 12544
rect 15252 12484 15256 12540
rect 15256 12484 15312 12540
rect 15312 12484 15316 12540
rect 15252 12480 15316 12484
rect 15332 12540 15396 12544
rect 15332 12484 15336 12540
rect 15336 12484 15392 12540
rect 15392 12484 15396 12540
rect 15332 12480 15396 12484
rect 15412 12540 15476 12544
rect 15412 12484 15416 12540
rect 15416 12484 15472 12540
rect 15472 12484 15476 12540
rect 15412 12480 15476 12484
rect 15492 12540 15556 12544
rect 15492 12484 15496 12540
rect 15496 12484 15552 12540
rect 15552 12484 15556 12540
rect 15492 12480 15556 12484
rect 18252 12540 18316 12544
rect 18252 12484 18256 12540
rect 18256 12484 18312 12540
rect 18312 12484 18316 12540
rect 18252 12480 18316 12484
rect 18332 12540 18396 12544
rect 18332 12484 18336 12540
rect 18336 12484 18392 12540
rect 18392 12484 18396 12540
rect 18332 12480 18396 12484
rect 18412 12540 18476 12544
rect 18412 12484 18416 12540
rect 18416 12484 18472 12540
rect 18472 12484 18476 12540
rect 18412 12480 18476 12484
rect 18492 12540 18556 12544
rect 18492 12484 18496 12540
rect 18496 12484 18552 12540
rect 18552 12484 18556 12540
rect 18492 12480 18556 12484
rect 21252 12540 21316 12544
rect 21252 12484 21256 12540
rect 21256 12484 21312 12540
rect 21312 12484 21316 12540
rect 21252 12480 21316 12484
rect 21332 12540 21396 12544
rect 21332 12484 21336 12540
rect 21336 12484 21392 12540
rect 21392 12484 21396 12540
rect 21332 12480 21396 12484
rect 21412 12540 21476 12544
rect 21412 12484 21416 12540
rect 21416 12484 21472 12540
rect 21472 12484 21476 12540
rect 21412 12480 21476 12484
rect 21492 12540 21556 12544
rect 21492 12484 21496 12540
rect 21496 12484 21552 12540
rect 21552 12484 21556 12540
rect 21492 12480 21556 12484
rect 24252 12540 24316 12544
rect 24252 12484 24256 12540
rect 24256 12484 24312 12540
rect 24312 12484 24316 12540
rect 24252 12480 24316 12484
rect 24332 12540 24396 12544
rect 24332 12484 24336 12540
rect 24336 12484 24392 12540
rect 24392 12484 24396 12540
rect 24332 12480 24396 12484
rect 24412 12540 24476 12544
rect 24412 12484 24416 12540
rect 24416 12484 24472 12540
rect 24472 12484 24476 12540
rect 24412 12480 24476 12484
rect 24492 12540 24556 12544
rect 24492 12484 24496 12540
rect 24496 12484 24552 12540
rect 24552 12484 24556 12540
rect 24492 12480 24556 12484
rect 27252 12540 27316 12544
rect 27252 12484 27256 12540
rect 27256 12484 27312 12540
rect 27312 12484 27316 12540
rect 27252 12480 27316 12484
rect 27332 12540 27396 12544
rect 27332 12484 27336 12540
rect 27336 12484 27392 12540
rect 27392 12484 27396 12540
rect 27332 12480 27396 12484
rect 27412 12540 27476 12544
rect 27412 12484 27416 12540
rect 27416 12484 27472 12540
rect 27472 12484 27476 12540
rect 27412 12480 27476 12484
rect 27492 12540 27556 12544
rect 27492 12484 27496 12540
rect 27496 12484 27552 12540
rect 27552 12484 27556 12540
rect 27492 12480 27556 12484
rect 1752 11996 1816 12000
rect 1752 11940 1756 11996
rect 1756 11940 1812 11996
rect 1812 11940 1816 11996
rect 1752 11936 1816 11940
rect 1832 11996 1896 12000
rect 1832 11940 1836 11996
rect 1836 11940 1892 11996
rect 1892 11940 1896 11996
rect 1832 11936 1896 11940
rect 1912 11996 1976 12000
rect 1912 11940 1916 11996
rect 1916 11940 1972 11996
rect 1972 11940 1976 11996
rect 1912 11936 1976 11940
rect 1992 11996 2056 12000
rect 1992 11940 1996 11996
rect 1996 11940 2052 11996
rect 2052 11940 2056 11996
rect 1992 11936 2056 11940
rect 4752 11996 4816 12000
rect 4752 11940 4756 11996
rect 4756 11940 4812 11996
rect 4812 11940 4816 11996
rect 4752 11936 4816 11940
rect 4832 11996 4896 12000
rect 4832 11940 4836 11996
rect 4836 11940 4892 11996
rect 4892 11940 4896 11996
rect 4832 11936 4896 11940
rect 4912 11996 4976 12000
rect 4912 11940 4916 11996
rect 4916 11940 4972 11996
rect 4972 11940 4976 11996
rect 4912 11936 4976 11940
rect 4992 11996 5056 12000
rect 4992 11940 4996 11996
rect 4996 11940 5052 11996
rect 5052 11940 5056 11996
rect 4992 11936 5056 11940
rect 7752 11996 7816 12000
rect 7752 11940 7756 11996
rect 7756 11940 7812 11996
rect 7812 11940 7816 11996
rect 7752 11936 7816 11940
rect 7832 11996 7896 12000
rect 7832 11940 7836 11996
rect 7836 11940 7892 11996
rect 7892 11940 7896 11996
rect 7832 11936 7896 11940
rect 7912 11996 7976 12000
rect 7912 11940 7916 11996
rect 7916 11940 7972 11996
rect 7972 11940 7976 11996
rect 7912 11936 7976 11940
rect 7992 11996 8056 12000
rect 7992 11940 7996 11996
rect 7996 11940 8052 11996
rect 8052 11940 8056 11996
rect 7992 11936 8056 11940
rect 10752 11996 10816 12000
rect 10752 11940 10756 11996
rect 10756 11940 10812 11996
rect 10812 11940 10816 11996
rect 10752 11936 10816 11940
rect 10832 11996 10896 12000
rect 10832 11940 10836 11996
rect 10836 11940 10892 11996
rect 10892 11940 10896 11996
rect 10832 11936 10896 11940
rect 10912 11996 10976 12000
rect 10912 11940 10916 11996
rect 10916 11940 10972 11996
rect 10972 11940 10976 11996
rect 10912 11936 10976 11940
rect 10992 11996 11056 12000
rect 10992 11940 10996 11996
rect 10996 11940 11052 11996
rect 11052 11940 11056 11996
rect 10992 11936 11056 11940
rect 13752 11996 13816 12000
rect 13752 11940 13756 11996
rect 13756 11940 13812 11996
rect 13812 11940 13816 11996
rect 13752 11936 13816 11940
rect 13832 11996 13896 12000
rect 13832 11940 13836 11996
rect 13836 11940 13892 11996
rect 13892 11940 13896 11996
rect 13832 11936 13896 11940
rect 13912 11996 13976 12000
rect 13912 11940 13916 11996
rect 13916 11940 13972 11996
rect 13972 11940 13976 11996
rect 13912 11936 13976 11940
rect 13992 11996 14056 12000
rect 13992 11940 13996 11996
rect 13996 11940 14052 11996
rect 14052 11940 14056 11996
rect 13992 11936 14056 11940
rect 16752 11996 16816 12000
rect 16752 11940 16756 11996
rect 16756 11940 16812 11996
rect 16812 11940 16816 11996
rect 16752 11936 16816 11940
rect 16832 11996 16896 12000
rect 16832 11940 16836 11996
rect 16836 11940 16892 11996
rect 16892 11940 16896 11996
rect 16832 11936 16896 11940
rect 16912 11996 16976 12000
rect 16912 11940 16916 11996
rect 16916 11940 16972 11996
rect 16972 11940 16976 11996
rect 16912 11936 16976 11940
rect 16992 11996 17056 12000
rect 16992 11940 16996 11996
rect 16996 11940 17052 11996
rect 17052 11940 17056 11996
rect 16992 11936 17056 11940
rect 19752 11996 19816 12000
rect 19752 11940 19756 11996
rect 19756 11940 19812 11996
rect 19812 11940 19816 11996
rect 19752 11936 19816 11940
rect 19832 11996 19896 12000
rect 19832 11940 19836 11996
rect 19836 11940 19892 11996
rect 19892 11940 19896 11996
rect 19832 11936 19896 11940
rect 19912 11996 19976 12000
rect 19912 11940 19916 11996
rect 19916 11940 19972 11996
rect 19972 11940 19976 11996
rect 19912 11936 19976 11940
rect 19992 11996 20056 12000
rect 19992 11940 19996 11996
rect 19996 11940 20052 11996
rect 20052 11940 20056 11996
rect 19992 11936 20056 11940
rect 22752 11996 22816 12000
rect 22752 11940 22756 11996
rect 22756 11940 22812 11996
rect 22812 11940 22816 11996
rect 22752 11936 22816 11940
rect 22832 11996 22896 12000
rect 22832 11940 22836 11996
rect 22836 11940 22892 11996
rect 22892 11940 22896 11996
rect 22832 11936 22896 11940
rect 22912 11996 22976 12000
rect 22912 11940 22916 11996
rect 22916 11940 22972 11996
rect 22972 11940 22976 11996
rect 22912 11936 22976 11940
rect 22992 11996 23056 12000
rect 22992 11940 22996 11996
rect 22996 11940 23052 11996
rect 23052 11940 23056 11996
rect 22992 11936 23056 11940
rect 25752 11996 25816 12000
rect 25752 11940 25756 11996
rect 25756 11940 25812 11996
rect 25812 11940 25816 11996
rect 25752 11936 25816 11940
rect 25832 11996 25896 12000
rect 25832 11940 25836 11996
rect 25836 11940 25892 11996
rect 25892 11940 25896 11996
rect 25832 11936 25896 11940
rect 25912 11996 25976 12000
rect 25912 11940 25916 11996
rect 25916 11940 25972 11996
rect 25972 11940 25976 11996
rect 25912 11936 25976 11940
rect 25992 11996 26056 12000
rect 25992 11940 25996 11996
rect 25996 11940 26052 11996
rect 26052 11940 26056 11996
rect 25992 11936 26056 11940
rect 3252 11452 3316 11456
rect 3252 11396 3256 11452
rect 3256 11396 3312 11452
rect 3312 11396 3316 11452
rect 3252 11392 3316 11396
rect 3332 11452 3396 11456
rect 3332 11396 3336 11452
rect 3336 11396 3392 11452
rect 3392 11396 3396 11452
rect 3332 11392 3396 11396
rect 3412 11452 3476 11456
rect 3412 11396 3416 11452
rect 3416 11396 3472 11452
rect 3472 11396 3476 11452
rect 3412 11392 3476 11396
rect 3492 11452 3556 11456
rect 3492 11396 3496 11452
rect 3496 11396 3552 11452
rect 3552 11396 3556 11452
rect 3492 11392 3556 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 6412 11452 6476 11456
rect 6412 11396 6416 11452
rect 6416 11396 6472 11452
rect 6472 11396 6476 11452
rect 6412 11392 6476 11396
rect 6492 11452 6556 11456
rect 6492 11396 6496 11452
rect 6496 11396 6552 11452
rect 6552 11396 6556 11452
rect 6492 11392 6556 11396
rect 9252 11452 9316 11456
rect 9252 11396 9256 11452
rect 9256 11396 9312 11452
rect 9312 11396 9316 11452
rect 9252 11392 9316 11396
rect 9332 11452 9396 11456
rect 9332 11396 9336 11452
rect 9336 11396 9392 11452
rect 9392 11396 9396 11452
rect 9332 11392 9396 11396
rect 9412 11452 9476 11456
rect 9412 11396 9416 11452
rect 9416 11396 9472 11452
rect 9472 11396 9476 11452
rect 9412 11392 9476 11396
rect 9492 11452 9556 11456
rect 9492 11396 9496 11452
rect 9496 11396 9552 11452
rect 9552 11396 9556 11452
rect 9492 11392 9556 11396
rect 12252 11452 12316 11456
rect 12252 11396 12256 11452
rect 12256 11396 12312 11452
rect 12312 11396 12316 11452
rect 12252 11392 12316 11396
rect 12332 11452 12396 11456
rect 12332 11396 12336 11452
rect 12336 11396 12392 11452
rect 12392 11396 12396 11452
rect 12332 11392 12396 11396
rect 12412 11452 12476 11456
rect 12412 11396 12416 11452
rect 12416 11396 12472 11452
rect 12472 11396 12476 11452
rect 12412 11392 12476 11396
rect 12492 11452 12556 11456
rect 12492 11396 12496 11452
rect 12496 11396 12552 11452
rect 12552 11396 12556 11452
rect 12492 11392 12556 11396
rect 15252 11452 15316 11456
rect 15252 11396 15256 11452
rect 15256 11396 15312 11452
rect 15312 11396 15316 11452
rect 15252 11392 15316 11396
rect 15332 11452 15396 11456
rect 15332 11396 15336 11452
rect 15336 11396 15392 11452
rect 15392 11396 15396 11452
rect 15332 11392 15396 11396
rect 15412 11452 15476 11456
rect 15412 11396 15416 11452
rect 15416 11396 15472 11452
rect 15472 11396 15476 11452
rect 15412 11392 15476 11396
rect 15492 11452 15556 11456
rect 15492 11396 15496 11452
rect 15496 11396 15552 11452
rect 15552 11396 15556 11452
rect 15492 11392 15556 11396
rect 18252 11452 18316 11456
rect 18252 11396 18256 11452
rect 18256 11396 18312 11452
rect 18312 11396 18316 11452
rect 18252 11392 18316 11396
rect 18332 11452 18396 11456
rect 18332 11396 18336 11452
rect 18336 11396 18392 11452
rect 18392 11396 18396 11452
rect 18332 11392 18396 11396
rect 18412 11452 18476 11456
rect 18412 11396 18416 11452
rect 18416 11396 18472 11452
rect 18472 11396 18476 11452
rect 18412 11392 18476 11396
rect 18492 11452 18556 11456
rect 18492 11396 18496 11452
rect 18496 11396 18552 11452
rect 18552 11396 18556 11452
rect 18492 11392 18556 11396
rect 21252 11452 21316 11456
rect 21252 11396 21256 11452
rect 21256 11396 21312 11452
rect 21312 11396 21316 11452
rect 21252 11392 21316 11396
rect 21332 11452 21396 11456
rect 21332 11396 21336 11452
rect 21336 11396 21392 11452
rect 21392 11396 21396 11452
rect 21332 11392 21396 11396
rect 21412 11452 21476 11456
rect 21412 11396 21416 11452
rect 21416 11396 21472 11452
rect 21472 11396 21476 11452
rect 21412 11392 21476 11396
rect 21492 11452 21556 11456
rect 21492 11396 21496 11452
rect 21496 11396 21552 11452
rect 21552 11396 21556 11452
rect 21492 11392 21556 11396
rect 24252 11452 24316 11456
rect 24252 11396 24256 11452
rect 24256 11396 24312 11452
rect 24312 11396 24316 11452
rect 24252 11392 24316 11396
rect 24332 11452 24396 11456
rect 24332 11396 24336 11452
rect 24336 11396 24392 11452
rect 24392 11396 24396 11452
rect 24332 11392 24396 11396
rect 24412 11452 24476 11456
rect 24412 11396 24416 11452
rect 24416 11396 24472 11452
rect 24472 11396 24476 11452
rect 24412 11392 24476 11396
rect 24492 11452 24556 11456
rect 24492 11396 24496 11452
rect 24496 11396 24552 11452
rect 24552 11396 24556 11452
rect 24492 11392 24556 11396
rect 27252 11452 27316 11456
rect 27252 11396 27256 11452
rect 27256 11396 27312 11452
rect 27312 11396 27316 11452
rect 27252 11392 27316 11396
rect 27332 11452 27396 11456
rect 27332 11396 27336 11452
rect 27336 11396 27392 11452
rect 27392 11396 27396 11452
rect 27332 11392 27396 11396
rect 27412 11452 27476 11456
rect 27412 11396 27416 11452
rect 27416 11396 27472 11452
rect 27472 11396 27476 11452
rect 27412 11392 27476 11396
rect 27492 11452 27556 11456
rect 27492 11396 27496 11452
rect 27496 11396 27552 11452
rect 27552 11396 27556 11452
rect 27492 11392 27556 11396
rect 1752 10908 1816 10912
rect 1752 10852 1756 10908
rect 1756 10852 1812 10908
rect 1812 10852 1816 10908
rect 1752 10848 1816 10852
rect 1832 10908 1896 10912
rect 1832 10852 1836 10908
rect 1836 10852 1892 10908
rect 1892 10852 1896 10908
rect 1832 10848 1896 10852
rect 1912 10908 1976 10912
rect 1912 10852 1916 10908
rect 1916 10852 1972 10908
rect 1972 10852 1976 10908
rect 1912 10848 1976 10852
rect 1992 10908 2056 10912
rect 1992 10852 1996 10908
rect 1996 10852 2052 10908
rect 2052 10852 2056 10908
rect 1992 10848 2056 10852
rect 4752 10908 4816 10912
rect 4752 10852 4756 10908
rect 4756 10852 4812 10908
rect 4812 10852 4816 10908
rect 4752 10848 4816 10852
rect 4832 10908 4896 10912
rect 4832 10852 4836 10908
rect 4836 10852 4892 10908
rect 4892 10852 4896 10908
rect 4832 10848 4896 10852
rect 4912 10908 4976 10912
rect 4912 10852 4916 10908
rect 4916 10852 4972 10908
rect 4972 10852 4976 10908
rect 4912 10848 4976 10852
rect 4992 10908 5056 10912
rect 4992 10852 4996 10908
rect 4996 10852 5052 10908
rect 5052 10852 5056 10908
rect 4992 10848 5056 10852
rect 7752 10908 7816 10912
rect 7752 10852 7756 10908
rect 7756 10852 7812 10908
rect 7812 10852 7816 10908
rect 7752 10848 7816 10852
rect 7832 10908 7896 10912
rect 7832 10852 7836 10908
rect 7836 10852 7892 10908
rect 7892 10852 7896 10908
rect 7832 10848 7896 10852
rect 7912 10908 7976 10912
rect 7912 10852 7916 10908
rect 7916 10852 7972 10908
rect 7972 10852 7976 10908
rect 7912 10848 7976 10852
rect 7992 10908 8056 10912
rect 7992 10852 7996 10908
rect 7996 10852 8052 10908
rect 8052 10852 8056 10908
rect 7992 10848 8056 10852
rect 10752 10908 10816 10912
rect 10752 10852 10756 10908
rect 10756 10852 10812 10908
rect 10812 10852 10816 10908
rect 10752 10848 10816 10852
rect 10832 10908 10896 10912
rect 10832 10852 10836 10908
rect 10836 10852 10892 10908
rect 10892 10852 10896 10908
rect 10832 10848 10896 10852
rect 10912 10908 10976 10912
rect 10912 10852 10916 10908
rect 10916 10852 10972 10908
rect 10972 10852 10976 10908
rect 10912 10848 10976 10852
rect 10992 10908 11056 10912
rect 10992 10852 10996 10908
rect 10996 10852 11052 10908
rect 11052 10852 11056 10908
rect 10992 10848 11056 10852
rect 13752 10908 13816 10912
rect 13752 10852 13756 10908
rect 13756 10852 13812 10908
rect 13812 10852 13816 10908
rect 13752 10848 13816 10852
rect 13832 10908 13896 10912
rect 13832 10852 13836 10908
rect 13836 10852 13892 10908
rect 13892 10852 13896 10908
rect 13832 10848 13896 10852
rect 13912 10908 13976 10912
rect 13912 10852 13916 10908
rect 13916 10852 13972 10908
rect 13972 10852 13976 10908
rect 13912 10848 13976 10852
rect 13992 10908 14056 10912
rect 13992 10852 13996 10908
rect 13996 10852 14052 10908
rect 14052 10852 14056 10908
rect 13992 10848 14056 10852
rect 16752 10908 16816 10912
rect 16752 10852 16756 10908
rect 16756 10852 16812 10908
rect 16812 10852 16816 10908
rect 16752 10848 16816 10852
rect 16832 10908 16896 10912
rect 16832 10852 16836 10908
rect 16836 10852 16892 10908
rect 16892 10852 16896 10908
rect 16832 10848 16896 10852
rect 16912 10908 16976 10912
rect 16912 10852 16916 10908
rect 16916 10852 16972 10908
rect 16972 10852 16976 10908
rect 16912 10848 16976 10852
rect 16992 10908 17056 10912
rect 16992 10852 16996 10908
rect 16996 10852 17052 10908
rect 17052 10852 17056 10908
rect 16992 10848 17056 10852
rect 19752 10908 19816 10912
rect 19752 10852 19756 10908
rect 19756 10852 19812 10908
rect 19812 10852 19816 10908
rect 19752 10848 19816 10852
rect 19832 10908 19896 10912
rect 19832 10852 19836 10908
rect 19836 10852 19892 10908
rect 19892 10852 19896 10908
rect 19832 10848 19896 10852
rect 19912 10908 19976 10912
rect 19912 10852 19916 10908
rect 19916 10852 19972 10908
rect 19972 10852 19976 10908
rect 19912 10848 19976 10852
rect 19992 10908 20056 10912
rect 19992 10852 19996 10908
rect 19996 10852 20052 10908
rect 20052 10852 20056 10908
rect 19992 10848 20056 10852
rect 22752 10908 22816 10912
rect 22752 10852 22756 10908
rect 22756 10852 22812 10908
rect 22812 10852 22816 10908
rect 22752 10848 22816 10852
rect 22832 10908 22896 10912
rect 22832 10852 22836 10908
rect 22836 10852 22892 10908
rect 22892 10852 22896 10908
rect 22832 10848 22896 10852
rect 22912 10908 22976 10912
rect 22912 10852 22916 10908
rect 22916 10852 22972 10908
rect 22972 10852 22976 10908
rect 22912 10848 22976 10852
rect 22992 10908 23056 10912
rect 22992 10852 22996 10908
rect 22996 10852 23052 10908
rect 23052 10852 23056 10908
rect 22992 10848 23056 10852
rect 25752 10908 25816 10912
rect 25752 10852 25756 10908
rect 25756 10852 25812 10908
rect 25812 10852 25816 10908
rect 25752 10848 25816 10852
rect 25832 10908 25896 10912
rect 25832 10852 25836 10908
rect 25836 10852 25892 10908
rect 25892 10852 25896 10908
rect 25832 10848 25896 10852
rect 25912 10908 25976 10912
rect 25912 10852 25916 10908
rect 25916 10852 25972 10908
rect 25972 10852 25976 10908
rect 25912 10848 25976 10852
rect 25992 10908 26056 10912
rect 25992 10852 25996 10908
rect 25996 10852 26052 10908
rect 26052 10852 26056 10908
rect 25992 10848 26056 10852
rect 3252 10364 3316 10368
rect 3252 10308 3256 10364
rect 3256 10308 3312 10364
rect 3312 10308 3316 10364
rect 3252 10304 3316 10308
rect 3332 10364 3396 10368
rect 3332 10308 3336 10364
rect 3336 10308 3392 10364
rect 3392 10308 3396 10364
rect 3332 10304 3396 10308
rect 3412 10364 3476 10368
rect 3412 10308 3416 10364
rect 3416 10308 3472 10364
rect 3472 10308 3476 10364
rect 3412 10304 3476 10308
rect 3492 10364 3556 10368
rect 3492 10308 3496 10364
rect 3496 10308 3552 10364
rect 3552 10308 3556 10364
rect 3492 10304 3556 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 6412 10364 6476 10368
rect 6412 10308 6416 10364
rect 6416 10308 6472 10364
rect 6472 10308 6476 10364
rect 6412 10304 6476 10308
rect 6492 10364 6556 10368
rect 6492 10308 6496 10364
rect 6496 10308 6552 10364
rect 6552 10308 6556 10364
rect 6492 10304 6556 10308
rect 9252 10364 9316 10368
rect 9252 10308 9256 10364
rect 9256 10308 9312 10364
rect 9312 10308 9316 10364
rect 9252 10304 9316 10308
rect 9332 10364 9396 10368
rect 9332 10308 9336 10364
rect 9336 10308 9392 10364
rect 9392 10308 9396 10364
rect 9332 10304 9396 10308
rect 9412 10364 9476 10368
rect 9412 10308 9416 10364
rect 9416 10308 9472 10364
rect 9472 10308 9476 10364
rect 9412 10304 9476 10308
rect 9492 10364 9556 10368
rect 9492 10308 9496 10364
rect 9496 10308 9552 10364
rect 9552 10308 9556 10364
rect 9492 10304 9556 10308
rect 12252 10364 12316 10368
rect 12252 10308 12256 10364
rect 12256 10308 12312 10364
rect 12312 10308 12316 10364
rect 12252 10304 12316 10308
rect 12332 10364 12396 10368
rect 12332 10308 12336 10364
rect 12336 10308 12392 10364
rect 12392 10308 12396 10364
rect 12332 10304 12396 10308
rect 12412 10364 12476 10368
rect 12412 10308 12416 10364
rect 12416 10308 12472 10364
rect 12472 10308 12476 10364
rect 12412 10304 12476 10308
rect 12492 10364 12556 10368
rect 12492 10308 12496 10364
rect 12496 10308 12552 10364
rect 12552 10308 12556 10364
rect 12492 10304 12556 10308
rect 15252 10364 15316 10368
rect 15252 10308 15256 10364
rect 15256 10308 15312 10364
rect 15312 10308 15316 10364
rect 15252 10304 15316 10308
rect 15332 10364 15396 10368
rect 15332 10308 15336 10364
rect 15336 10308 15392 10364
rect 15392 10308 15396 10364
rect 15332 10304 15396 10308
rect 15412 10364 15476 10368
rect 15412 10308 15416 10364
rect 15416 10308 15472 10364
rect 15472 10308 15476 10364
rect 15412 10304 15476 10308
rect 15492 10364 15556 10368
rect 15492 10308 15496 10364
rect 15496 10308 15552 10364
rect 15552 10308 15556 10364
rect 15492 10304 15556 10308
rect 18252 10364 18316 10368
rect 18252 10308 18256 10364
rect 18256 10308 18312 10364
rect 18312 10308 18316 10364
rect 18252 10304 18316 10308
rect 18332 10364 18396 10368
rect 18332 10308 18336 10364
rect 18336 10308 18392 10364
rect 18392 10308 18396 10364
rect 18332 10304 18396 10308
rect 18412 10364 18476 10368
rect 18412 10308 18416 10364
rect 18416 10308 18472 10364
rect 18472 10308 18476 10364
rect 18412 10304 18476 10308
rect 18492 10364 18556 10368
rect 18492 10308 18496 10364
rect 18496 10308 18552 10364
rect 18552 10308 18556 10364
rect 18492 10304 18556 10308
rect 21252 10364 21316 10368
rect 21252 10308 21256 10364
rect 21256 10308 21312 10364
rect 21312 10308 21316 10364
rect 21252 10304 21316 10308
rect 21332 10364 21396 10368
rect 21332 10308 21336 10364
rect 21336 10308 21392 10364
rect 21392 10308 21396 10364
rect 21332 10304 21396 10308
rect 21412 10364 21476 10368
rect 21412 10308 21416 10364
rect 21416 10308 21472 10364
rect 21472 10308 21476 10364
rect 21412 10304 21476 10308
rect 21492 10364 21556 10368
rect 21492 10308 21496 10364
rect 21496 10308 21552 10364
rect 21552 10308 21556 10364
rect 21492 10304 21556 10308
rect 24252 10364 24316 10368
rect 24252 10308 24256 10364
rect 24256 10308 24312 10364
rect 24312 10308 24316 10364
rect 24252 10304 24316 10308
rect 24332 10364 24396 10368
rect 24332 10308 24336 10364
rect 24336 10308 24392 10364
rect 24392 10308 24396 10364
rect 24332 10304 24396 10308
rect 24412 10364 24476 10368
rect 24412 10308 24416 10364
rect 24416 10308 24472 10364
rect 24472 10308 24476 10364
rect 24412 10304 24476 10308
rect 24492 10364 24556 10368
rect 24492 10308 24496 10364
rect 24496 10308 24552 10364
rect 24552 10308 24556 10364
rect 24492 10304 24556 10308
rect 27252 10364 27316 10368
rect 27252 10308 27256 10364
rect 27256 10308 27312 10364
rect 27312 10308 27316 10364
rect 27252 10304 27316 10308
rect 27332 10364 27396 10368
rect 27332 10308 27336 10364
rect 27336 10308 27392 10364
rect 27392 10308 27396 10364
rect 27332 10304 27396 10308
rect 27412 10364 27476 10368
rect 27412 10308 27416 10364
rect 27416 10308 27472 10364
rect 27472 10308 27476 10364
rect 27412 10304 27476 10308
rect 27492 10364 27556 10368
rect 27492 10308 27496 10364
rect 27496 10308 27552 10364
rect 27552 10308 27556 10364
rect 27492 10304 27556 10308
rect 1752 9820 1816 9824
rect 1752 9764 1756 9820
rect 1756 9764 1812 9820
rect 1812 9764 1816 9820
rect 1752 9760 1816 9764
rect 1832 9820 1896 9824
rect 1832 9764 1836 9820
rect 1836 9764 1892 9820
rect 1892 9764 1896 9820
rect 1832 9760 1896 9764
rect 1912 9820 1976 9824
rect 1912 9764 1916 9820
rect 1916 9764 1972 9820
rect 1972 9764 1976 9820
rect 1912 9760 1976 9764
rect 1992 9820 2056 9824
rect 1992 9764 1996 9820
rect 1996 9764 2052 9820
rect 2052 9764 2056 9820
rect 1992 9760 2056 9764
rect 4752 9820 4816 9824
rect 4752 9764 4756 9820
rect 4756 9764 4812 9820
rect 4812 9764 4816 9820
rect 4752 9760 4816 9764
rect 4832 9820 4896 9824
rect 4832 9764 4836 9820
rect 4836 9764 4892 9820
rect 4892 9764 4896 9820
rect 4832 9760 4896 9764
rect 4912 9820 4976 9824
rect 4912 9764 4916 9820
rect 4916 9764 4972 9820
rect 4972 9764 4976 9820
rect 4912 9760 4976 9764
rect 4992 9820 5056 9824
rect 4992 9764 4996 9820
rect 4996 9764 5052 9820
rect 5052 9764 5056 9820
rect 4992 9760 5056 9764
rect 7752 9820 7816 9824
rect 7752 9764 7756 9820
rect 7756 9764 7812 9820
rect 7812 9764 7816 9820
rect 7752 9760 7816 9764
rect 7832 9820 7896 9824
rect 7832 9764 7836 9820
rect 7836 9764 7892 9820
rect 7892 9764 7896 9820
rect 7832 9760 7896 9764
rect 7912 9820 7976 9824
rect 7912 9764 7916 9820
rect 7916 9764 7972 9820
rect 7972 9764 7976 9820
rect 7912 9760 7976 9764
rect 7992 9820 8056 9824
rect 7992 9764 7996 9820
rect 7996 9764 8052 9820
rect 8052 9764 8056 9820
rect 7992 9760 8056 9764
rect 10752 9820 10816 9824
rect 10752 9764 10756 9820
rect 10756 9764 10812 9820
rect 10812 9764 10816 9820
rect 10752 9760 10816 9764
rect 10832 9820 10896 9824
rect 10832 9764 10836 9820
rect 10836 9764 10892 9820
rect 10892 9764 10896 9820
rect 10832 9760 10896 9764
rect 10912 9820 10976 9824
rect 10912 9764 10916 9820
rect 10916 9764 10972 9820
rect 10972 9764 10976 9820
rect 10912 9760 10976 9764
rect 10992 9820 11056 9824
rect 10992 9764 10996 9820
rect 10996 9764 11052 9820
rect 11052 9764 11056 9820
rect 10992 9760 11056 9764
rect 13752 9820 13816 9824
rect 13752 9764 13756 9820
rect 13756 9764 13812 9820
rect 13812 9764 13816 9820
rect 13752 9760 13816 9764
rect 13832 9820 13896 9824
rect 13832 9764 13836 9820
rect 13836 9764 13892 9820
rect 13892 9764 13896 9820
rect 13832 9760 13896 9764
rect 13912 9820 13976 9824
rect 13912 9764 13916 9820
rect 13916 9764 13972 9820
rect 13972 9764 13976 9820
rect 13912 9760 13976 9764
rect 13992 9820 14056 9824
rect 13992 9764 13996 9820
rect 13996 9764 14052 9820
rect 14052 9764 14056 9820
rect 13992 9760 14056 9764
rect 16752 9820 16816 9824
rect 16752 9764 16756 9820
rect 16756 9764 16812 9820
rect 16812 9764 16816 9820
rect 16752 9760 16816 9764
rect 16832 9820 16896 9824
rect 16832 9764 16836 9820
rect 16836 9764 16892 9820
rect 16892 9764 16896 9820
rect 16832 9760 16896 9764
rect 16912 9820 16976 9824
rect 16912 9764 16916 9820
rect 16916 9764 16972 9820
rect 16972 9764 16976 9820
rect 16912 9760 16976 9764
rect 16992 9820 17056 9824
rect 16992 9764 16996 9820
rect 16996 9764 17052 9820
rect 17052 9764 17056 9820
rect 16992 9760 17056 9764
rect 19752 9820 19816 9824
rect 19752 9764 19756 9820
rect 19756 9764 19812 9820
rect 19812 9764 19816 9820
rect 19752 9760 19816 9764
rect 19832 9820 19896 9824
rect 19832 9764 19836 9820
rect 19836 9764 19892 9820
rect 19892 9764 19896 9820
rect 19832 9760 19896 9764
rect 19912 9820 19976 9824
rect 19912 9764 19916 9820
rect 19916 9764 19972 9820
rect 19972 9764 19976 9820
rect 19912 9760 19976 9764
rect 19992 9820 20056 9824
rect 19992 9764 19996 9820
rect 19996 9764 20052 9820
rect 20052 9764 20056 9820
rect 19992 9760 20056 9764
rect 22752 9820 22816 9824
rect 22752 9764 22756 9820
rect 22756 9764 22812 9820
rect 22812 9764 22816 9820
rect 22752 9760 22816 9764
rect 22832 9820 22896 9824
rect 22832 9764 22836 9820
rect 22836 9764 22892 9820
rect 22892 9764 22896 9820
rect 22832 9760 22896 9764
rect 22912 9820 22976 9824
rect 22912 9764 22916 9820
rect 22916 9764 22972 9820
rect 22972 9764 22976 9820
rect 22912 9760 22976 9764
rect 22992 9820 23056 9824
rect 22992 9764 22996 9820
rect 22996 9764 23052 9820
rect 23052 9764 23056 9820
rect 22992 9760 23056 9764
rect 25752 9820 25816 9824
rect 25752 9764 25756 9820
rect 25756 9764 25812 9820
rect 25812 9764 25816 9820
rect 25752 9760 25816 9764
rect 25832 9820 25896 9824
rect 25832 9764 25836 9820
rect 25836 9764 25892 9820
rect 25892 9764 25896 9820
rect 25832 9760 25896 9764
rect 25912 9820 25976 9824
rect 25912 9764 25916 9820
rect 25916 9764 25972 9820
rect 25972 9764 25976 9820
rect 25912 9760 25976 9764
rect 25992 9820 26056 9824
rect 25992 9764 25996 9820
rect 25996 9764 26052 9820
rect 26052 9764 26056 9820
rect 25992 9760 26056 9764
rect 3252 9276 3316 9280
rect 3252 9220 3256 9276
rect 3256 9220 3312 9276
rect 3312 9220 3316 9276
rect 3252 9216 3316 9220
rect 3332 9276 3396 9280
rect 3332 9220 3336 9276
rect 3336 9220 3392 9276
rect 3392 9220 3396 9276
rect 3332 9216 3396 9220
rect 3412 9276 3476 9280
rect 3412 9220 3416 9276
rect 3416 9220 3472 9276
rect 3472 9220 3476 9276
rect 3412 9216 3476 9220
rect 3492 9276 3556 9280
rect 3492 9220 3496 9276
rect 3496 9220 3552 9276
rect 3552 9220 3556 9276
rect 3492 9216 3556 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 6412 9276 6476 9280
rect 6412 9220 6416 9276
rect 6416 9220 6472 9276
rect 6472 9220 6476 9276
rect 6412 9216 6476 9220
rect 6492 9276 6556 9280
rect 6492 9220 6496 9276
rect 6496 9220 6552 9276
rect 6552 9220 6556 9276
rect 6492 9216 6556 9220
rect 9252 9276 9316 9280
rect 9252 9220 9256 9276
rect 9256 9220 9312 9276
rect 9312 9220 9316 9276
rect 9252 9216 9316 9220
rect 9332 9276 9396 9280
rect 9332 9220 9336 9276
rect 9336 9220 9392 9276
rect 9392 9220 9396 9276
rect 9332 9216 9396 9220
rect 9412 9276 9476 9280
rect 9412 9220 9416 9276
rect 9416 9220 9472 9276
rect 9472 9220 9476 9276
rect 9412 9216 9476 9220
rect 9492 9276 9556 9280
rect 9492 9220 9496 9276
rect 9496 9220 9552 9276
rect 9552 9220 9556 9276
rect 9492 9216 9556 9220
rect 12252 9276 12316 9280
rect 12252 9220 12256 9276
rect 12256 9220 12312 9276
rect 12312 9220 12316 9276
rect 12252 9216 12316 9220
rect 12332 9276 12396 9280
rect 12332 9220 12336 9276
rect 12336 9220 12392 9276
rect 12392 9220 12396 9276
rect 12332 9216 12396 9220
rect 12412 9276 12476 9280
rect 12412 9220 12416 9276
rect 12416 9220 12472 9276
rect 12472 9220 12476 9276
rect 12412 9216 12476 9220
rect 12492 9276 12556 9280
rect 12492 9220 12496 9276
rect 12496 9220 12552 9276
rect 12552 9220 12556 9276
rect 12492 9216 12556 9220
rect 15252 9276 15316 9280
rect 15252 9220 15256 9276
rect 15256 9220 15312 9276
rect 15312 9220 15316 9276
rect 15252 9216 15316 9220
rect 15332 9276 15396 9280
rect 15332 9220 15336 9276
rect 15336 9220 15392 9276
rect 15392 9220 15396 9276
rect 15332 9216 15396 9220
rect 15412 9276 15476 9280
rect 15412 9220 15416 9276
rect 15416 9220 15472 9276
rect 15472 9220 15476 9276
rect 15412 9216 15476 9220
rect 15492 9276 15556 9280
rect 15492 9220 15496 9276
rect 15496 9220 15552 9276
rect 15552 9220 15556 9276
rect 15492 9216 15556 9220
rect 18252 9276 18316 9280
rect 18252 9220 18256 9276
rect 18256 9220 18312 9276
rect 18312 9220 18316 9276
rect 18252 9216 18316 9220
rect 18332 9276 18396 9280
rect 18332 9220 18336 9276
rect 18336 9220 18392 9276
rect 18392 9220 18396 9276
rect 18332 9216 18396 9220
rect 18412 9276 18476 9280
rect 18412 9220 18416 9276
rect 18416 9220 18472 9276
rect 18472 9220 18476 9276
rect 18412 9216 18476 9220
rect 18492 9276 18556 9280
rect 18492 9220 18496 9276
rect 18496 9220 18552 9276
rect 18552 9220 18556 9276
rect 18492 9216 18556 9220
rect 21252 9276 21316 9280
rect 21252 9220 21256 9276
rect 21256 9220 21312 9276
rect 21312 9220 21316 9276
rect 21252 9216 21316 9220
rect 21332 9276 21396 9280
rect 21332 9220 21336 9276
rect 21336 9220 21392 9276
rect 21392 9220 21396 9276
rect 21332 9216 21396 9220
rect 21412 9276 21476 9280
rect 21412 9220 21416 9276
rect 21416 9220 21472 9276
rect 21472 9220 21476 9276
rect 21412 9216 21476 9220
rect 21492 9276 21556 9280
rect 21492 9220 21496 9276
rect 21496 9220 21552 9276
rect 21552 9220 21556 9276
rect 21492 9216 21556 9220
rect 24252 9276 24316 9280
rect 24252 9220 24256 9276
rect 24256 9220 24312 9276
rect 24312 9220 24316 9276
rect 24252 9216 24316 9220
rect 24332 9276 24396 9280
rect 24332 9220 24336 9276
rect 24336 9220 24392 9276
rect 24392 9220 24396 9276
rect 24332 9216 24396 9220
rect 24412 9276 24476 9280
rect 24412 9220 24416 9276
rect 24416 9220 24472 9276
rect 24472 9220 24476 9276
rect 24412 9216 24476 9220
rect 24492 9276 24556 9280
rect 24492 9220 24496 9276
rect 24496 9220 24552 9276
rect 24552 9220 24556 9276
rect 24492 9216 24556 9220
rect 27252 9276 27316 9280
rect 27252 9220 27256 9276
rect 27256 9220 27312 9276
rect 27312 9220 27316 9276
rect 27252 9216 27316 9220
rect 27332 9276 27396 9280
rect 27332 9220 27336 9276
rect 27336 9220 27392 9276
rect 27392 9220 27396 9276
rect 27332 9216 27396 9220
rect 27412 9276 27476 9280
rect 27412 9220 27416 9276
rect 27416 9220 27472 9276
rect 27472 9220 27476 9276
rect 27412 9216 27476 9220
rect 27492 9276 27556 9280
rect 27492 9220 27496 9276
rect 27496 9220 27552 9276
rect 27552 9220 27556 9276
rect 27492 9216 27556 9220
rect 1752 8732 1816 8736
rect 1752 8676 1756 8732
rect 1756 8676 1812 8732
rect 1812 8676 1816 8732
rect 1752 8672 1816 8676
rect 1832 8732 1896 8736
rect 1832 8676 1836 8732
rect 1836 8676 1892 8732
rect 1892 8676 1896 8732
rect 1832 8672 1896 8676
rect 1912 8732 1976 8736
rect 1912 8676 1916 8732
rect 1916 8676 1972 8732
rect 1972 8676 1976 8732
rect 1912 8672 1976 8676
rect 1992 8732 2056 8736
rect 1992 8676 1996 8732
rect 1996 8676 2052 8732
rect 2052 8676 2056 8732
rect 1992 8672 2056 8676
rect 4752 8732 4816 8736
rect 4752 8676 4756 8732
rect 4756 8676 4812 8732
rect 4812 8676 4816 8732
rect 4752 8672 4816 8676
rect 4832 8732 4896 8736
rect 4832 8676 4836 8732
rect 4836 8676 4892 8732
rect 4892 8676 4896 8732
rect 4832 8672 4896 8676
rect 4912 8732 4976 8736
rect 4912 8676 4916 8732
rect 4916 8676 4972 8732
rect 4972 8676 4976 8732
rect 4912 8672 4976 8676
rect 4992 8732 5056 8736
rect 4992 8676 4996 8732
rect 4996 8676 5052 8732
rect 5052 8676 5056 8732
rect 4992 8672 5056 8676
rect 7752 8732 7816 8736
rect 7752 8676 7756 8732
rect 7756 8676 7812 8732
rect 7812 8676 7816 8732
rect 7752 8672 7816 8676
rect 7832 8732 7896 8736
rect 7832 8676 7836 8732
rect 7836 8676 7892 8732
rect 7892 8676 7896 8732
rect 7832 8672 7896 8676
rect 7912 8732 7976 8736
rect 7912 8676 7916 8732
rect 7916 8676 7972 8732
rect 7972 8676 7976 8732
rect 7912 8672 7976 8676
rect 7992 8732 8056 8736
rect 7992 8676 7996 8732
rect 7996 8676 8052 8732
rect 8052 8676 8056 8732
rect 7992 8672 8056 8676
rect 10752 8732 10816 8736
rect 10752 8676 10756 8732
rect 10756 8676 10812 8732
rect 10812 8676 10816 8732
rect 10752 8672 10816 8676
rect 10832 8732 10896 8736
rect 10832 8676 10836 8732
rect 10836 8676 10892 8732
rect 10892 8676 10896 8732
rect 10832 8672 10896 8676
rect 10912 8732 10976 8736
rect 10912 8676 10916 8732
rect 10916 8676 10972 8732
rect 10972 8676 10976 8732
rect 10912 8672 10976 8676
rect 10992 8732 11056 8736
rect 10992 8676 10996 8732
rect 10996 8676 11052 8732
rect 11052 8676 11056 8732
rect 10992 8672 11056 8676
rect 13752 8732 13816 8736
rect 13752 8676 13756 8732
rect 13756 8676 13812 8732
rect 13812 8676 13816 8732
rect 13752 8672 13816 8676
rect 13832 8732 13896 8736
rect 13832 8676 13836 8732
rect 13836 8676 13892 8732
rect 13892 8676 13896 8732
rect 13832 8672 13896 8676
rect 13912 8732 13976 8736
rect 13912 8676 13916 8732
rect 13916 8676 13972 8732
rect 13972 8676 13976 8732
rect 13912 8672 13976 8676
rect 13992 8732 14056 8736
rect 13992 8676 13996 8732
rect 13996 8676 14052 8732
rect 14052 8676 14056 8732
rect 13992 8672 14056 8676
rect 16752 8732 16816 8736
rect 16752 8676 16756 8732
rect 16756 8676 16812 8732
rect 16812 8676 16816 8732
rect 16752 8672 16816 8676
rect 16832 8732 16896 8736
rect 16832 8676 16836 8732
rect 16836 8676 16892 8732
rect 16892 8676 16896 8732
rect 16832 8672 16896 8676
rect 16912 8732 16976 8736
rect 16912 8676 16916 8732
rect 16916 8676 16972 8732
rect 16972 8676 16976 8732
rect 16912 8672 16976 8676
rect 16992 8732 17056 8736
rect 16992 8676 16996 8732
rect 16996 8676 17052 8732
rect 17052 8676 17056 8732
rect 16992 8672 17056 8676
rect 19752 8732 19816 8736
rect 19752 8676 19756 8732
rect 19756 8676 19812 8732
rect 19812 8676 19816 8732
rect 19752 8672 19816 8676
rect 19832 8732 19896 8736
rect 19832 8676 19836 8732
rect 19836 8676 19892 8732
rect 19892 8676 19896 8732
rect 19832 8672 19896 8676
rect 19912 8732 19976 8736
rect 19912 8676 19916 8732
rect 19916 8676 19972 8732
rect 19972 8676 19976 8732
rect 19912 8672 19976 8676
rect 19992 8732 20056 8736
rect 19992 8676 19996 8732
rect 19996 8676 20052 8732
rect 20052 8676 20056 8732
rect 19992 8672 20056 8676
rect 22752 8732 22816 8736
rect 22752 8676 22756 8732
rect 22756 8676 22812 8732
rect 22812 8676 22816 8732
rect 22752 8672 22816 8676
rect 22832 8732 22896 8736
rect 22832 8676 22836 8732
rect 22836 8676 22892 8732
rect 22892 8676 22896 8732
rect 22832 8672 22896 8676
rect 22912 8732 22976 8736
rect 22912 8676 22916 8732
rect 22916 8676 22972 8732
rect 22972 8676 22976 8732
rect 22912 8672 22976 8676
rect 22992 8732 23056 8736
rect 22992 8676 22996 8732
rect 22996 8676 23052 8732
rect 23052 8676 23056 8732
rect 22992 8672 23056 8676
rect 25752 8732 25816 8736
rect 25752 8676 25756 8732
rect 25756 8676 25812 8732
rect 25812 8676 25816 8732
rect 25752 8672 25816 8676
rect 25832 8732 25896 8736
rect 25832 8676 25836 8732
rect 25836 8676 25892 8732
rect 25892 8676 25896 8732
rect 25832 8672 25896 8676
rect 25912 8732 25976 8736
rect 25912 8676 25916 8732
rect 25916 8676 25972 8732
rect 25972 8676 25976 8732
rect 25912 8672 25976 8676
rect 25992 8732 26056 8736
rect 25992 8676 25996 8732
rect 25996 8676 26052 8732
rect 26052 8676 26056 8732
rect 25992 8672 26056 8676
rect 3252 8188 3316 8192
rect 3252 8132 3256 8188
rect 3256 8132 3312 8188
rect 3312 8132 3316 8188
rect 3252 8128 3316 8132
rect 3332 8188 3396 8192
rect 3332 8132 3336 8188
rect 3336 8132 3392 8188
rect 3392 8132 3396 8188
rect 3332 8128 3396 8132
rect 3412 8188 3476 8192
rect 3412 8132 3416 8188
rect 3416 8132 3472 8188
rect 3472 8132 3476 8188
rect 3412 8128 3476 8132
rect 3492 8188 3556 8192
rect 3492 8132 3496 8188
rect 3496 8132 3552 8188
rect 3552 8132 3556 8188
rect 3492 8128 3556 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 6412 8188 6476 8192
rect 6412 8132 6416 8188
rect 6416 8132 6472 8188
rect 6472 8132 6476 8188
rect 6412 8128 6476 8132
rect 6492 8188 6556 8192
rect 6492 8132 6496 8188
rect 6496 8132 6552 8188
rect 6552 8132 6556 8188
rect 6492 8128 6556 8132
rect 9252 8188 9316 8192
rect 9252 8132 9256 8188
rect 9256 8132 9312 8188
rect 9312 8132 9316 8188
rect 9252 8128 9316 8132
rect 9332 8188 9396 8192
rect 9332 8132 9336 8188
rect 9336 8132 9392 8188
rect 9392 8132 9396 8188
rect 9332 8128 9396 8132
rect 9412 8188 9476 8192
rect 9412 8132 9416 8188
rect 9416 8132 9472 8188
rect 9472 8132 9476 8188
rect 9412 8128 9476 8132
rect 9492 8188 9556 8192
rect 9492 8132 9496 8188
rect 9496 8132 9552 8188
rect 9552 8132 9556 8188
rect 9492 8128 9556 8132
rect 12252 8188 12316 8192
rect 12252 8132 12256 8188
rect 12256 8132 12312 8188
rect 12312 8132 12316 8188
rect 12252 8128 12316 8132
rect 12332 8188 12396 8192
rect 12332 8132 12336 8188
rect 12336 8132 12392 8188
rect 12392 8132 12396 8188
rect 12332 8128 12396 8132
rect 12412 8188 12476 8192
rect 12412 8132 12416 8188
rect 12416 8132 12472 8188
rect 12472 8132 12476 8188
rect 12412 8128 12476 8132
rect 12492 8188 12556 8192
rect 12492 8132 12496 8188
rect 12496 8132 12552 8188
rect 12552 8132 12556 8188
rect 12492 8128 12556 8132
rect 15252 8188 15316 8192
rect 15252 8132 15256 8188
rect 15256 8132 15312 8188
rect 15312 8132 15316 8188
rect 15252 8128 15316 8132
rect 15332 8188 15396 8192
rect 15332 8132 15336 8188
rect 15336 8132 15392 8188
rect 15392 8132 15396 8188
rect 15332 8128 15396 8132
rect 15412 8188 15476 8192
rect 15412 8132 15416 8188
rect 15416 8132 15472 8188
rect 15472 8132 15476 8188
rect 15412 8128 15476 8132
rect 15492 8188 15556 8192
rect 15492 8132 15496 8188
rect 15496 8132 15552 8188
rect 15552 8132 15556 8188
rect 15492 8128 15556 8132
rect 18252 8188 18316 8192
rect 18252 8132 18256 8188
rect 18256 8132 18312 8188
rect 18312 8132 18316 8188
rect 18252 8128 18316 8132
rect 18332 8188 18396 8192
rect 18332 8132 18336 8188
rect 18336 8132 18392 8188
rect 18392 8132 18396 8188
rect 18332 8128 18396 8132
rect 18412 8188 18476 8192
rect 18412 8132 18416 8188
rect 18416 8132 18472 8188
rect 18472 8132 18476 8188
rect 18412 8128 18476 8132
rect 18492 8188 18556 8192
rect 18492 8132 18496 8188
rect 18496 8132 18552 8188
rect 18552 8132 18556 8188
rect 18492 8128 18556 8132
rect 21252 8188 21316 8192
rect 21252 8132 21256 8188
rect 21256 8132 21312 8188
rect 21312 8132 21316 8188
rect 21252 8128 21316 8132
rect 21332 8188 21396 8192
rect 21332 8132 21336 8188
rect 21336 8132 21392 8188
rect 21392 8132 21396 8188
rect 21332 8128 21396 8132
rect 21412 8188 21476 8192
rect 21412 8132 21416 8188
rect 21416 8132 21472 8188
rect 21472 8132 21476 8188
rect 21412 8128 21476 8132
rect 21492 8188 21556 8192
rect 21492 8132 21496 8188
rect 21496 8132 21552 8188
rect 21552 8132 21556 8188
rect 21492 8128 21556 8132
rect 24252 8188 24316 8192
rect 24252 8132 24256 8188
rect 24256 8132 24312 8188
rect 24312 8132 24316 8188
rect 24252 8128 24316 8132
rect 24332 8188 24396 8192
rect 24332 8132 24336 8188
rect 24336 8132 24392 8188
rect 24392 8132 24396 8188
rect 24332 8128 24396 8132
rect 24412 8188 24476 8192
rect 24412 8132 24416 8188
rect 24416 8132 24472 8188
rect 24472 8132 24476 8188
rect 24412 8128 24476 8132
rect 24492 8188 24556 8192
rect 24492 8132 24496 8188
rect 24496 8132 24552 8188
rect 24552 8132 24556 8188
rect 24492 8128 24556 8132
rect 27252 8188 27316 8192
rect 27252 8132 27256 8188
rect 27256 8132 27312 8188
rect 27312 8132 27316 8188
rect 27252 8128 27316 8132
rect 27332 8188 27396 8192
rect 27332 8132 27336 8188
rect 27336 8132 27392 8188
rect 27392 8132 27396 8188
rect 27332 8128 27396 8132
rect 27412 8188 27476 8192
rect 27412 8132 27416 8188
rect 27416 8132 27472 8188
rect 27472 8132 27476 8188
rect 27412 8128 27476 8132
rect 27492 8188 27556 8192
rect 27492 8132 27496 8188
rect 27496 8132 27552 8188
rect 27552 8132 27556 8188
rect 27492 8128 27556 8132
rect 1752 7644 1816 7648
rect 1752 7588 1756 7644
rect 1756 7588 1812 7644
rect 1812 7588 1816 7644
rect 1752 7584 1816 7588
rect 1832 7644 1896 7648
rect 1832 7588 1836 7644
rect 1836 7588 1892 7644
rect 1892 7588 1896 7644
rect 1832 7584 1896 7588
rect 1912 7644 1976 7648
rect 1912 7588 1916 7644
rect 1916 7588 1972 7644
rect 1972 7588 1976 7644
rect 1912 7584 1976 7588
rect 1992 7644 2056 7648
rect 1992 7588 1996 7644
rect 1996 7588 2052 7644
rect 2052 7588 2056 7644
rect 1992 7584 2056 7588
rect 4752 7644 4816 7648
rect 4752 7588 4756 7644
rect 4756 7588 4812 7644
rect 4812 7588 4816 7644
rect 4752 7584 4816 7588
rect 4832 7644 4896 7648
rect 4832 7588 4836 7644
rect 4836 7588 4892 7644
rect 4892 7588 4896 7644
rect 4832 7584 4896 7588
rect 4912 7644 4976 7648
rect 4912 7588 4916 7644
rect 4916 7588 4972 7644
rect 4972 7588 4976 7644
rect 4912 7584 4976 7588
rect 4992 7644 5056 7648
rect 4992 7588 4996 7644
rect 4996 7588 5052 7644
rect 5052 7588 5056 7644
rect 4992 7584 5056 7588
rect 7752 7644 7816 7648
rect 7752 7588 7756 7644
rect 7756 7588 7812 7644
rect 7812 7588 7816 7644
rect 7752 7584 7816 7588
rect 7832 7644 7896 7648
rect 7832 7588 7836 7644
rect 7836 7588 7892 7644
rect 7892 7588 7896 7644
rect 7832 7584 7896 7588
rect 7912 7644 7976 7648
rect 7912 7588 7916 7644
rect 7916 7588 7972 7644
rect 7972 7588 7976 7644
rect 7912 7584 7976 7588
rect 7992 7644 8056 7648
rect 7992 7588 7996 7644
rect 7996 7588 8052 7644
rect 8052 7588 8056 7644
rect 7992 7584 8056 7588
rect 10752 7644 10816 7648
rect 10752 7588 10756 7644
rect 10756 7588 10812 7644
rect 10812 7588 10816 7644
rect 10752 7584 10816 7588
rect 10832 7644 10896 7648
rect 10832 7588 10836 7644
rect 10836 7588 10892 7644
rect 10892 7588 10896 7644
rect 10832 7584 10896 7588
rect 10912 7644 10976 7648
rect 10912 7588 10916 7644
rect 10916 7588 10972 7644
rect 10972 7588 10976 7644
rect 10912 7584 10976 7588
rect 10992 7644 11056 7648
rect 10992 7588 10996 7644
rect 10996 7588 11052 7644
rect 11052 7588 11056 7644
rect 10992 7584 11056 7588
rect 13752 7644 13816 7648
rect 13752 7588 13756 7644
rect 13756 7588 13812 7644
rect 13812 7588 13816 7644
rect 13752 7584 13816 7588
rect 13832 7644 13896 7648
rect 13832 7588 13836 7644
rect 13836 7588 13892 7644
rect 13892 7588 13896 7644
rect 13832 7584 13896 7588
rect 13912 7644 13976 7648
rect 13912 7588 13916 7644
rect 13916 7588 13972 7644
rect 13972 7588 13976 7644
rect 13912 7584 13976 7588
rect 13992 7644 14056 7648
rect 13992 7588 13996 7644
rect 13996 7588 14052 7644
rect 14052 7588 14056 7644
rect 13992 7584 14056 7588
rect 16752 7644 16816 7648
rect 16752 7588 16756 7644
rect 16756 7588 16812 7644
rect 16812 7588 16816 7644
rect 16752 7584 16816 7588
rect 16832 7644 16896 7648
rect 16832 7588 16836 7644
rect 16836 7588 16892 7644
rect 16892 7588 16896 7644
rect 16832 7584 16896 7588
rect 16912 7644 16976 7648
rect 16912 7588 16916 7644
rect 16916 7588 16972 7644
rect 16972 7588 16976 7644
rect 16912 7584 16976 7588
rect 16992 7644 17056 7648
rect 16992 7588 16996 7644
rect 16996 7588 17052 7644
rect 17052 7588 17056 7644
rect 16992 7584 17056 7588
rect 19752 7644 19816 7648
rect 19752 7588 19756 7644
rect 19756 7588 19812 7644
rect 19812 7588 19816 7644
rect 19752 7584 19816 7588
rect 19832 7644 19896 7648
rect 19832 7588 19836 7644
rect 19836 7588 19892 7644
rect 19892 7588 19896 7644
rect 19832 7584 19896 7588
rect 19912 7644 19976 7648
rect 19912 7588 19916 7644
rect 19916 7588 19972 7644
rect 19972 7588 19976 7644
rect 19912 7584 19976 7588
rect 19992 7644 20056 7648
rect 19992 7588 19996 7644
rect 19996 7588 20052 7644
rect 20052 7588 20056 7644
rect 19992 7584 20056 7588
rect 22752 7644 22816 7648
rect 22752 7588 22756 7644
rect 22756 7588 22812 7644
rect 22812 7588 22816 7644
rect 22752 7584 22816 7588
rect 22832 7644 22896 7648
rect 22832 7588 22836 7644
rect 22836 7588 22892 7644
rect 22892 7588 22896 7644
rect 22832 7584 22896 7588
rect 22912 7644 22976 7648
rect 22912 7588 22916 7644
rect 22916 7588 22972 7644
rect 22972 7588 22976 7644
rect 22912 7584 22976 7588
rect 22992 7644 23056 7648
rect 22992 7588 22996 7644
rect 22996 7588 23052 7644
rect 23052 7588 23056 7644
rect 22992 7584 23056 7588
rect 25752 7644 25816 7648
rect 25752 7588 25756 7644
rect 25756 7588 25812 7644
rect 25812 7588 25816 7644
rect 25752 7584 25816 7588
rect 25832 7644 25896 7648
rect 25832 7588 25836 7644
rect 25836 7588 25892 7644
rect 25892 7588 25896 7644
rect 25832 7584 25896 7588
rect 25912 7644 25976 7648
rect 25912 7588 25916 7644
rect 25916 7588 25972 7644
rect 25972 7588 25976 7644
rect 25912 7584 25976 7588
rect 25992 7644 26056 7648
rect 25992 7588 25996 7644
rect 25996 7588 26052 7644
rect 26052 7588 26056 7644
rect 25992 7584 26056 7588
rect 3252 7100 3316 7104
rect 3252 7044 3256 7100
rect 3256 7044 3312 7100
rect 3312 7044 3316 7100
rect 3252 7040 3316 7044
rect 3332 7100 3396 7104
rect 3332 7044 3336 7100
rect 3336 7044 3392 7100
rect 3392 7044 3396 7100
rect 3332 7040 3396 7044
rect 3412 7100 3476 7104
rect 3412 7044 3416 7100
rect 3416 7044 3472 7100
rect 3472 7044 3476 7100
rect 3412 7040 3476 7044
rect 3492 7100 3556 7104
rect 3492 7044 3496 7100
rect 3496 7044 3552 7100
rect 3552 7044 3556 7100
rect 3492 7040 3556 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 6412 7100 6476 7104
rect 6412 7044 6416 7100
rect 6416 7044 6472 7100
rect 6472 7044 6476 7100
rect 6412 7040 6476 7044
rect 6492 7100 6556 7104
rect 6492 7044 6496 7100
rect 6496 7044 6552 7100
rect 6552 7044 6556 7100
rect 6492 7040 6556 7044
rect 9252 7100 9316 7104
rect 9252 7044 9256 7100
rect 9256 7044 9312 7100
rect 9312 7044 9316 7100
rect 9252 7040 9316 7044
rect 9332 7100 9396 7104
rect 9332 7044 9336 7100
rect 9336 7044 9392 7100
rect 9392 7044 9396 7100
rect 9332 7040 9396 7044
rect 9412 7100 9476 7104
rect 9412 7044 9416 7100
rect 9416 7044 9472 7100
rect 9472 7044 9476 7100
rect 9412 7040 9476 7044
rect 9492 7100 9556 7104
rect 9492 7044 9496 7100
rect 9496 7044 9552 7100
rect 9552 7044 9556 7100
rect 9492 7040 9556 7044
rect 12252 7100 12316 7104
rect 12252 7044 12256 7100
rect 12256 7044 12312 7100
rect 12312 7044 12316 7100
rect 12252 7040 12316 7044
rect 12332 7100 12396 7104
rect 12332 7044 12336 7100
rect 12336 7044 12392 7100
rect 12392 7044 12396 7100
rect 12332 7040 12396 7044
rect 12412 7100 12476 7104
rect 12412 7044 12416 7100
rect 12416 7044 12472 7100
rect 12472 7044 12476 7100
rect 12412 7040 12476 7044
rect 12492 7100 12556 7104
rect 12492 7044 12496 7100
rect 12496 7044 12552 7100
rect 12552 7044 12556 7100
rect 12492 7040 12556 7044
rect 15252 7100 15316 7104
rect 15252 7044 15256 7100
rect 15256 7044 15312 7100
rect 15312 7044 15316 7100
rect 15252 7040 15316 7044
rect 15332 7100 15396 7104
rect 15332 7044 15336 7100
rect 15336 7044 15392 7100
rect 15392 7044 15396 7100
rect 15332 7040 15396 7044
rect 15412 7100 15476 7104
rect 15412 7044 15416 7100
rect 15416 7044 15472 7100
rect 15472 7044 15476 7100
rect 15412 7040 15476 7044
rect 15492 7100 15556 7104
rect 15492 7044 15496 7100
rect 15496 7044 15552 7100
rect 15552 7044 15556 7100
rect 15492 7040 15556 7044
rect 18252 7100 18316 7104
rect 18252 7044 18256 7100
rect 18256 7044 18312 7100
rect 18312 7044 18316 7100
rect 18252 7040 18316 7044
rect 18332 7100 18396 7104
rect 18332 7044 18336 7100
rect 18336 7044 18392 7100
rect 18392 7044 18396 7100
rect 18332 7040 18396 7044
rect 18412 7100 18476 7104
rect 18412 7044 18416 7100
rect 18416 7044 18472 7100
rect 18472 7044 18476 7100
rect 18412 7040 18476 7044
rect 18492 7100 18556 7104
rect 18492 7044 18496 7100
rect 18496 7044 18552 7100
rect 18552 7044 18556 7100
rect 18492 7040 18556 7044
rect 21252 7100 21316 7104
rect 21252 7044 21256 7100
rect 21256 7044 21312 7100
rect 21312 7044 21316 7100
rect 21252 7040 21316 7044
rect 21332 7100 21396 7104
rect 21332 7044 21336 7100
rect 21336 7044 21392 7100
rect 21392 7044 21396 7100
rect 21332 7040 21396 7044
rect 21412 7100 21476 7104
rect 21412 7044 21416 7100
rect 21416 7044 21472 7100
rect 21472 7044 21476 7100
rect 21412 7040 21476 7044
rect 21492 7100 21556 7104
rect 21492 7044 21496 7100
rect 21496 7044 21552 7100
rect 21552 7044 21556 7100
rect 21492 7040 21556 7044
rect 24252 7100 24316 7104
rect 24252 7044 24256 7100
rect 24256 7044 24312 7100
rect 24312 7044 24316 7100
rect 24252 7040 24316 7044
rect 24332 7100 24396 7104
rect 24332 7044 24336 7100
rect 24336 7044 24392 7100
rect 24392 7044 24396 7100
rect 24332 7040 24396 7044
rect 24412 7100 24476 7104
rect 24412 7044 24416 7100
rect 24416 7044 24472 7100
rect 24472 7044 24476 7100
rect 24412 7040 24476 7044
rect 24492 7100 24556 7104
rect 24492 7044 24496 7100
rect 24496 7044 24552 7100
rect 24552 7044 24556 7100
rect 24492 7040 24556 7044
rect 27252 7100 27316 7104
rect 27252 7044 27256 7100
rect 27256 7044 27312 7100
rect 27312 7044 27316 7100
rect 27252 7040 27316 7044
rect 27332 7100 27396 7104
rect 27332 7044 27336 7100
rect 27336 7044 27392 7100
rect 27392 7044 27396 7100
rect 27332 7040 27396 7044
rect 27412 7100 27476 7104
rect 27412 7044 27416 7100
rect 27416 7044 27472 7100
rect 27472 7044 27476 7100
rect 27412 7040 27476 7044
rect 27492 7100 27556 7104
rect 27492 7044 27496 7100
rect 27496 7044 27552 7100
rect 27552 7044 27556 7100
rect 27492 7040 27556 7044
rect 1752 6556 1816 6560
rect 1752 6500 1756 6556
rect 1756 6500 1812 6556
rect 1812 6500 1816 6556
rect 1752 6496 1816 6500
rect 1832 6556 1896 6560
rect 1832 6500 1836 6556
rect 1836 6500 1892 6556
rect 1892 6500 1896 6556
rect 1832 6496 1896 6500
rect 1912 6556 1976 6560
rect 1912 6500 1916 6556
rect 1916 6500 1972 6556
rect 1972 6500 1976 6556
rect 1912 6496 1976 6500
rect 1992 6556 2056 6560
rect 1992 6500 1996 6556
rect 1996 6500 2052 6556
rect 2052 6500 2056 6556
rect 1992 6496 2056 6500
rect 4752 6556 4816 6560
rect 4752 6500 4756 6556
rect 4756 6500 4812 6556
rect 4812 6500 4816 6556
rect 4752 6496 4816 6500
rect 4832 6556 4896 6560
rect 4832 6500 4836 6556
rect 4836 6500 4892 6556
rect 4892 6500 4896 6556
rect 4832 6496 4896 6500
rect 4912 6556 4976 6560
rect 4912 6500 4916 6556
rect 4916 6500 4972 6556
rect 4972 6500 4976 6556
rect 4912 6496 4976 6500
rect 4992 6556 5056 6560
rect 4992 6500 4996 6556
rect 4996 6500 5052 6556
rect 5052 6500 5056 6556
rect 4992 6496 5056 6500
rect 7752 6556 7816 6560
rect 7752 6500 7756 6556
rect 7756 6500 7812 6556
rect 7812 6500 7816 6556
rect 7752 6496 7816 6500
rect 7832 6556 7896 6560
rect 7832 6500 7836 6556
rect 7836 6500 7892 6556
rect 7892 6500 7896 6556
rect 7832 6496 7896 6500
rect 7912 6556 7976 6560
rect 7912 6500 7916 6556
rect 7916 6500 7972 6556
rect 7972 6500 7976 6556
rect 7912 6496 7976 6500
rect 7992 6556 8056 6560
rect 7992 6500 7996 6556
rect 7996 6500 8052 6556
rect 8052 6500 8056 6556
rect 7992 6496 8056 6500
rect 10752 6556 10816 6560
rect 10752 6500 10756 6556
rect 10756 6500 10812 6556
rect 10812 6500 10816 6556
rect 10752 6496 10816 6500
rect 10832 6556 10896 6560
rect 10832 6500 10836 6556
rect 10836 6500 10892 6556
rect 10892 6500 10896 6556
rect 10832 6496 10896 6500
rect 10912 6556 10976 6560
rect 10912 6500 10916 6556
rect 10916 6500 10972 6556
rect 10972 6500 10976 6556
rect 10912 6496 10976 6500
rect 10992 6556 11056 6560
rect 10992 6500 10996 6556
rect 10996 6500 11052 6556
rect 11052 6500 11056 6556
rect 10992 6496 11056 6500
rect 13752 6556 13816 6560
rect 13752 6500 13756 6556
rect 13756 6500 13812 6556
rect 13812 6500 13816 6556
rect 13752 6496 13816 6500
rect 13832 6556 13896 6560
rect 13832 6500 13836 6556
rect 13836 6500 13892 6556
rect 13892 6500 13896 6556
rect 13832 6496 13896 6500
rect 13912 6556 13976 6560
rect 13912 6500 13916 6556
rect 13916 6500 13972 6556
rect 13972 6500 13976 6556
rect 13912 6496 13976 6500
rect 13992 6556 14056 6560
rect 13992 6500 13996 6556
rect 13996 6500 14052 6556
rect 14052 6500 14056 6556
rect 13992 6496 14056 6500
rect 16752 6556 16816 6560
rect 16752 6500 16756 6556
rect 16756 6500 16812 6556
rect 16812 6500 16816 6556
rect 16752 6496 16816 6500
rect 16832 6556 16896 6560
rect 16832 6500 16836 6556
rect 16836 6500 16892 6556
rect 16892 6500 16896 6556
rect 16832 6496 16896 6500
rect 16912 6556 16976 6560
rect 16912 6500 16916 6556
rect 16916 6500 16972 6556
rect 16972 6500 16976 6556
rect 16912 6496 16976 6500
rect 16992 6556 17056 6560
rect 16992 6500 16996 6556
rect 16996 6500 17052 6556
rect 17052 6500 17056 6556
rect 16992 6496 17056 6500
rect 19752 6556 19816 6560
rect 19752 6500 19756 6556
rect 19756 6500 19812 6556
rect 19812 6500 19816 6556
rect 19752 6496 19816 6500
rect 19832 6556 19896 6560
rect 19832 6500 19836 6556
rect 19836 6500 19892 6556
rect 19892 6500 19896 6556
rect 19832 6496 19896 6500
rect 19912 6556 19976 6560
rect 19912 6500 19916 6556
rect 19916 6500 19972 6556
rect 19972 6500 19976 6556
rect 19912 6496 19976 6500
rect 19992 6556 20056 6560
rect 19992 6500 19996 6556
rect 19996 6500 20052 6556
rect 20052 6500 20056 6556
rect 19992 6496 20056 6500
rect 22752 6556 22816 6560
rect 22752 6500 22756 6556
rect 22756 6500 22812 6556
rect 22812 6500 22816 6556
rect 22752 6496 22816 6500
rect 22832 6556 22896 6560
rect 22832 6500 22836 6556
rect 22836 6500 22892 6556
rect 22892 6500 22896 6556
rect 22832 6496 22896 6500
rect 22912 6556 22976 6560
rect 22912 6500 22916 6556
rect 22916 6500 22972 6556
rect 22972 6500 22976 6556
rect 22912 6496 22976 6500
rect 22992 6556 23056 6560
rect 22992 6500 22996 6556
rect 22996 6500 23052 6556
rect 23052 6500 23056 6556
rect 22992 6496 23056 6500
rect 25752 6556 25816 6560
rect 25752 6500 25756 6556
rect 25756 6500 25812 6556
rect 25812 6500 25816 6556
rect 25752 6496 25816 6500
rect 25832 6556 25896 6560
rect 25832 6500 25836 6556
rect 25836 6500 25892 6556
rect 25892 6500 25896 6556
rect 25832 6496 25896 6500
rect 25912 6556 25976 6560
rect 25912 6500 25916 6556
rect 25916 6500 25972 6556
rect 25972 6500 25976 6556
rect 25912 6496 25976 6500
rect 25992 6556 26056 6560
rect 25992 6500 25996 6556
rect 25996 6500 26052 6556
rect 26052 6500 26056 6556
rect 25992 6496 26056 6500
rect 3252 6012 3316 6016
rect 3252 5956 3256 6012
rect 3256 5956 3312 6012
rect 3312 5956 3316 6012
rect 3252 5952 3316 5956
rect 3332 6012 3396 6016
rect 3332 5956 3336 6012
rect 3336 5956 3392 6012
rect 3392 5956 3396 6012
rect 3332 5952 3396 5956
rect 3412 6012 3476 6016
rect 3412 5956 3416 6012
rect 3416 5956 3472 6012
rect 3472 5956 3476 6012
rect 3412 5952 3476 5956
rect 3492 6012 3556 6016
rect 3492 5956 3496 6012
rect 3496 5956 3552 6012
rect 3552 5956 3556 6012
rect 3492 5952 3556 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 6412 6012 6476 6016
rect 6412 5956 6416 6012
rect 6416 5956 6472 6012
rect 6472 5956 6476 6012
rect 6412 5952 6476 5956
rect 6492 6012 6556 6016
rect 6492 5956 6496 6012
rect 6496 5956 6552 6012
rect 6552 5956 6556 6012
rect 6492 5952 6556 5956
rect 9252 6012 9316 6016
rect 9252 5956 9256 6012
rect 9256 5956 9312 6012
rect 9312 5956 9316 6012
rect 9252 5952 9316 5956
rect 9332 6012 9396 6016
rect 9332 5956 9336 6012
rect 9336 5956 9392 6012
rect 9392 5956 9396 6012
rect 9332 5952 9396 5956
rect 9412 6012 9476 6016
rect 9412 5956 9416 6012
rect 9416 5956 9472 6012
rect 9472 5956 9476 6012
rect 9412 5952 9476 5956
rect 9492 6012 9556 6016
rect 9492 5956 9496 6012
rect 9496 5956 9552 6012
rect 9552 5956 9556 6012
rect 9492 5952 9556 5956
rect 12252 6012 12316 6016
rect 12252 5956 12256 6012
rect 12256 5956 12312 6012
rect 12312 5956 12316 6012
rect 12252 5952 12316 5956
rect 12332 6012 12396 6016
rect 12332 5956 12336 6012
rect 12336 5956 12392 6012
rect 12392 5956 12396 6012
rect 12332 5952 12396 5956
rect 12412 6012 12476 6016
rect 12412 5956 12416 6012
rect 12416 5956 12472 6012
rect 12472 5956 12476 6012
rect 12412 5952 12476 5956
rect 12492 6012 12556 6016
rect 12492 5956 12496 6012
rect 12496 5956 12552 6012
rect 12552 5956 12556 6012
rect 12492 5952 12556 5956
rect 15252 6012 15316 6016
rect 15252 5956 15256 6012
rect 15256 5956 15312 6012
rect 15312 5956 15316 6012
rect 15252 5952 15316 5956
rect 15332 6012 15396 6016
rect 15332 5956 15336 6012
rect 15336 5956 15392 6012
rect 15392 5956 15396 6012
rect 15332 5952 15396 5956
rect 15412 6012 15476 6016
rect 15412 5956 15416 6012
rect 15416 5956 15472 6012
rect 15472 5956 15476 6012
rect 15412 5952 15476 5956
rect 15492 6012 15556 6016
rect 15492 5956 15496 6012
rect 15496 5956 15552 6012
rect 15552 5956 15556 6012
rect 15492 5952 15556 5956
rect 18252 6012 18316 6016
rect 18252 5956 18256 6012
rect 18256 5956 18312 6012
rect 18312 5956 18316 6012
rect 18252 5952 18316 5956
rect 18332 6012 18396 6016
rect 18332 5956 18336 6012
rect 18336 5956 18392 6012
rect 18392 5956 18396 6012
rect 18332 5952 18396 5956
rect 18412 6012 18476 6016
rect 18412 5956 18416 6012
rect 18416 5956 18472 6012
rect 18472 5956 18476 6012
rect 18412 5952 18476 5956
rect 18492 6012 18556 6016
rect 18492 5956 18496 6012
rect 18496 5956 18552 6012
rect 18552 5956 18556 6012
rect 18492 5952 18556 5956
rect 21252 6012 21316 6016
rect 21252 5956 21256 6012
rect 21256 5956 21312 6012
rect 21312 5956 21316 6012
rect 21252 5952 21316 5956
rect 21332 6012 21396 6016
rect 21332 5956 21336 6012
rect 21336 5956 21392 6012
rect 21392 5956 21396 6012
rect 21332 5952 21396 5956
rect 21412 6012 21476 6016
rect 21412 5956 21416 6012
rect 21416 5956 21472 6012
rect 21472 5956 21476 6012
rect 21412 5952 21476 5956
rect 21492 6012 21556 6016
rect 21492 5956 21496 6012
rect 21496 5956 21552 6012
rect 21552 5956 21556 6012
rect 21492 5952 21556 5956
rect 24252 6012 24316 6016
rect 24252 5956 24256 6012
rect 24256 5956 24312 6012
rect 24312 5956 24316 6012
rect 24252 5952 24316 5956
rect 24332 6012 24396 6016
rect 24332 5956 24336 6012
rect 24336 5956 24392 6012
rect 24392 5956 24396 6012
rect 24332 5952 24396 5956
rect 24412 6012 24476 6016
rect 24412 5956 24416 6012
rect 24416 5956 24472 6012
rect 24472 5956 24476 6012
rect 24412 5952 24476 5956
rect 24492 6012 24556 6016
rect 24492 5956 24496 6012
rect 24496 5956 24552 6012
rect 24552 5956 24556 6012
rect 24492 5952 24556 5956
rect 27252 6012 27316 6016
rect 27252 5956 27256 6012
rect 27256 5956 27312 6012
rect 27312 5956 27316 6012
rect 27252 5952 27316 5956
rect 27332 6012 27396 6016
rect 27332 5956 27336 6012
rect 27336 5956 27392 6012
rect 27392 5956 27396 6012
rect 27332 5952 27396 5956
rect 27412 6012 27476 6016
rect 27412 5956 27416 6012
rect 27416 5956 27472 6012
rect 27472 5956 27476 6012
rect 27412 5952 27476 5956
rect 27492 6012 27556 6016
rect 27492 5956 27496 6012
rect 27496 5956 27552 6012
rect 27552 5956 27556 6012
rect 27492 5952 27556 5956
rect 1752 5468 1816 5472
rect 1752 5412 1756 5468
rect 1756 5412 1812 5468
rect 1812 5412 1816 5468
rect 1752 5408 1816 5412
rect 1832 5468 1896 5472
rect 1832 5412 1836 5468
rect 1836 5412 1892 5468
rect 1892 5412 1896 5468
rect 1832 5408 1896 5412
rect 1912 5468 1976 5472
rect 1912 5412 1916 5468
rect 1916 5412 1972 5468
rect 1972 5412 1976 5468
rect 1912 5408 1976 5412
rect 1992 5468 2056 5472
rect 1992 5412 1996 5468
rect 1996 5412 2052 5468
rect 2052 5412 2056 5468
rect 1992 5408 2056 5412
rect 4752 5468 4816 5472
rect 4752 5412 4756 5468
rect 4756 5412 4812 5468
rect 4812 5412 4816 5468
rect 4752 5408 4816 5412
rect 4832 5468 4896 5472
rect 4832 5412 4836 5468
rect 4836 5412 4892 5468
rect 4892 5412 4896 5468
rect 4832 5408 4896 5412
rect 4912 5468 4976 5472
rect 4912 5412 4916 5468
rect 4916 5412 4972 5468
rect 4972 5412 4976 5468
rect 4912 5408 4976 5412
rect 4992 5468 5056 5472
rect 4992 5412 4996 5468
rect 4996 5412 5052 5468
rect 5052 5412 5056 5468
rect 4992 5408 5056 5412
rect 7752 5468 7816 5472
rect 7752 5412 7756 5468
rect 7756 5412 7812 5468
rect 7812 5412 7816 5468
rect 7752 5408 7816 5412
rect 7832 5468 7896 5472
rect 7832 5412 7836 5468
rect 7836 5412 7892 5468
rect 7892 5412 7896 5468
rect 7832 5408 7896 5412
rect 7912 5468 7976 5472
rect 7912 5412 7916 5468
rect 7916 5412 7972 5468
rect 7972 5412 7976 5468
rect 7912 5408 7976 5412
rect 7992 5468 8056 5472
rect 7992 5412 7996 5468
rect 7996 5412 8052 5468
rect 8052 5412 8056 5468
rect 7992 5408 8056 5412
rect 10752 5468 10816 5472
rect 10752 5412 10756 5468
rect 10756 5412 10812 5468
rect 10812 5412 10816 5468
rect 10752 5408 10816 5412
rect 10832 5468 10896 5472
rect 10832 5412 10836 5468
rect 10836 5412 10892 5468
rect 10892 5412 10896 5468
rect 10832 5408 10896 5412
rect 10912 5468 10976 5472
rect 10912 5412 10916 5468
rect 10916 5412 10972 5468
rect 10972 5412 10976 5468
rect 10912 5408 10976 5412
rect 10992 5468 11056 5472
rect 10992 5412 10996 5468
rect 10996 5412 11052 5468
rect 11052 5412 11056 5468
rect 10992 5408 11056 5412
rect 13752 5468 13816 5472
rect 13752 5412 13756 5468
rect 13756 5412 13812 5468
rect 13812 5412 13816 5468
rect 13752 5408 13816 5412
rect 13832 5468 13896 5472
rect 13832 5412 13836 5468
rect 13836 5412 13892 5468
rect 13892 5412 13896 5468
rect 13832 5408 13896 5412
rect 13912 5468 13976 5472
rect 13912 5412 13916 5468
rect 13916 5412 13972 5468
rect 13972 5412 13976 5468
rect 13912 5408 13976 5412
rect 13992 5468 14056 5472
rect 13992 5412 13996 5468
rect 13996 5412 14052 5468
rect 14052 5412 14056 5468
rect 13992 5408 14056 5412
rect 16752 5468 16816 5472
rect 16752 5412 16756 5468
rect 16756 5412 16812 5468
rect 16812 5412 16816 5468
rect 16752 5408 16816 5412
rect 16832 5468 16896 5472
rect 16832 5412 16836 5468
rect 16836 5412 16892 5468
rect 16892 5412 16896 5468
rect 16832 5408 16896 5412
rect 16912 5468 16976 5472
rect 16912 5412 16916 5468
rect 16916 5412 16972 5468
rect 16972 5412 16976 5468
rect 16912 5408 16976 5412
rect 16992 5468 17056 5472
rect 16992 5412 16996 5468
rect 16996 5412 17052 5468
rect 17052 5412 17056 5468
rect 16992 5408 17056 5412
rect 19752 5468 19816 5472
rect 19752 5412 19756 5468
rect 19756 5412 19812 5468
rect 19812 5412 19816 5468
rect 19752 5408 19816 5412
rect 19832 5468 19896 5472
rect 19832 5412 19836 5468
rect 19836 5412 19892 5468
rect 19892 5412 19896 5468
rect 19832 5408 19896 5412
rect 19912 5468 19976 5472
rect 19912 5412 19916 5468
rect 19916 5412 19972 5468
rect 19972 5412 19976 5468
rect 19912 5408 19976 5412
rect 19992 5468 20056 5472
rect 19992 5412 19996 5468
rect 19996 5412 20052 5468
rect 20052 5412 20056 5468
rect 19992 5408 20056 5412
rect 22752 5468 22816 5472
rect 22752 5412 22756 5468
rect 22756 5412 22812 5468
rect 22812 5412 22816 5468
rect 22752 5408 22816 5412
rect 22832 5468 22896 5472
rect 22832 5412 22836 5468
rect 22836 5412 22892 5468
rect 22892 5412 22896 5468
rect 22832 5408 22896 5412
rect 22912 5468 22976 5472
rect 22912 5412 22916 5468
rect 22916 5412 22972 5468
rect 22972 5412 22976 5468
rect 22912 5408 22976 5412
rect 22992 5468 23056 5472
rect 22992 5412 22996 5468
rect 22996 5412 23052 5468
rect 23052 5412 23056 5468
rect 22992 5408 23056 5412
rect 25752 5468 25816 5472
rect 25752 5412 25756 5468
rect 25756 5412 25812 5468
rect 25812 5412 25816 5468
rect 25752 5408 25816 5412
rect 25832 5468 25896 5472
rect 25832 5412 25836 5468
rect 25836 5412 25892 5468
rect 25892 5412 25896 5468
rect 25832 5408 25896 5412
rect 25912 5468 25976 5472
rect 25912 5412 25916 5468
rect 25916 5412 25972 5468
rect 25972 5412 25976 5468
rect 25912 5408 25976 5412
rect 25992 5468 26056 5472
rect 25992 5412 25996 5468
rect 25996 5412 26052 5468
rect 26052 5412 26056 5468
rect 25992 5408 26056 5412
rect 3252 4924 3316 4928
rect 3252 4868 3256 4924
rect 3256 4868 3312 4924
rect 3312 4868 3316 4924
rect 3252 4864 3316 4868
rect 3332 4924 3396 4928
rect 3332 4868 3336 4924
rect 3336 4868 3392 4924
rect 3392 4868 3396 4924
rect 3332 4864 3396 4868
rect 3412 4924 3476 4928
rect 3412 4868 3416 4924
rect 3416 4868 3472 4924
rect 3472 4868 3476 4924
rect 3412 4864 3476 4868
rect 3492 4924 3556 4928
rect 3492 4868 3496 4924
rect 3496 4868 3552 4924
rect 3552 4868 3556 4924
rect 3492 4864 3556 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 6412 4924 6476 4928
rect 6412 4868 6416 4924
rect 6416 4868 6472 4924
rect 6472 4868 6476 4924
rect 6412 4864 6476 4868
rect 6492 4924 6556 4928
rect 6492 4868 6496 4924
rect 6496 4868 6552 4924
rect 6552 4868 6556 4924
rect 6492 4864 6556 4868
rect 9252 4924 9316 4928
rect 9252 4868 9256 4924
rect 9256 4868 9312 4924
rect 9312 4868 9316 4924
rect 9252 4864 9316 4868
rect 9332 4924 9396 4928
rect 9332 4868 9336 4924
rect 9336 4868 9392 4924
rect 9392 4868 9396 4924
rect 9332 4864 9396 4868
rect 9412 4924 9476 4928
rect 9412 4868 9416 4924
rect 9416 4868 9472 4924
rect 9472 4868 9476 4924
rect 9412 4864 9476 4868
rect 9492 4924 9556 4928
rect 9492 4868 9496 4924
rect 9496 4868 9552 4924
rect 9552 4868 9556 4924
rect 9492 4864 9556 4868
rect 12252 4924 12316 4928
rect 12252 4868 12256 4924
rect 12256 4868 12312 4924
rect 12312 4868 12316 4924
rect 12252 4864 12316 4868
rect 12332 4924 12396 4928
rect 12332 4868 12336 4924
rect 12336 4868 12392 4924
rect 12392 4868 12396 4924
rect 12332 4864 12396 4868
rect 12412 4924 12476 4928
rect 12412 4868 12416 4924
rect 12416 4868 12472 4924
rect 12472 4868 12476 4924
rect 12412 4864 12476 4868
rect 12492 4924 12556 4928
rect 12492 4868 12496 4924
rect 12496 4868 12552 4924
rect 12552 4868 12556 4924
rect 12492 4864 12556 4868
rect 15252 4924 15316 4928
rect 15252 4868 15256 4924
rect 15256 4868 15312 4924
rect 15312 4868 15316 4924
rect 15252 4864 15316 4868
rect 15332 4924 15396 4928
rect 15332 4868 15336 4924
rect 15336 4868 15392 4924
rect 15392 4868 15396 4924
rect 15332 4864 15396 4868
rect 15412 4924 15476 4928
rect 15412 4868 15416 4924
rect 15416 4868 15472 4924
rect 15472 4868 15476 4924
rect 15412 4864 15476 4868
rect 15492 4924 15556 4928
rect 15492 4868 15496 4924
rect 15496 4868 15552 4924
rect 15552 4868 15556 4924
rect 15492 4864 15556 4868
rect 18252 4924 18316 4928
rect 18252 4868 18256 4924
rect 18256 4868 18312 4924
rect 18312 4868 18316 4924
rect 18252 4864 18316 4868
rect 18332 4924 18396 4928
rect 18332 4868 18336 4924
rect 18336 4868 18392 4924
rect 18392 4868 18396 4924
rect 18332 4864 18396 4868
rect 18412 4924 18476 4928
rect 18412 4868 18416 4924
rect 18416 4868 18472 4924
rect 18472 4868 18476 4924
rect 18412 4864 18476 4868
rect 18492 4924 18556 4928
rect 18492 4868 18496 4924
rect 18496 4868 18552 4924
rect 18552 4868 18556 4924
rect 18492 4864 18556 4868
rect 21252 4924 21316 4928
rect 21252 4868 21256 4924
rect 21256 4868 21312 4924
rect 21312 4868 21316 4924
rect 21252 4864 21316 4868
rect 21332 4924 21396 4928
rect 21332 4868 21336 4924
rect 21336 4868 21392 4924
rect 21392 4868 21396 4924
rect 21332 4864 21396 4868
rect 21412 4924 21476 4928
rect 21412 4868 21416 4924
rect 21416 4868 21472 4924
rect 21472 4868 21476 4924
rect 21412 4864 21476 4868
rect 21492 4924 21556 4928
rect 21492 4868 21496 4924
rect 21496 4868 21552 4924
rect 21552 4868 21556 4924
rect 21492 4864 21556 4868
rect 24252 4924 24316 4928
rect 24252 4868 24256 4924
rect 24256 4868 24312 4924
rect 24312 4868 24316 4924
rect 24252 4864 24316 4868
rect 24332 4924 24396 4928
rect 24332 4868 24336 4924
rect 24336 4868 24392 4924
rect 24392 4868 24396 4924
rect 24332 4864 24396 4868
rect 24412 4924 24476 4928
rect 24412 4868 24416 4924
rect 24416 4868 24472 4924
rect 24472 4868 24476 4924
rect 24412 4864 24476 4868
rect 24492 4924 24556 4928
rect 24492 4868 24496 4924
rect 24496 4868 24552 4924
rect 24552 4868 24556 4924
rect 24492 4864 24556 4868
rect 27252 4924 27316 4928
rect 27252 4868 27256 4924
rect 27256 4868 27312 4924
rect 27312 4868 27316 4924
rect 27252 4864 27316 4868
rect 27332 4924 27396 4928
rect 27332 4868 27336 4924
rect 27336 4868 27392 4924
rect 27392 4868 27396 4924
rect 27332 4864 27396 4868
rect 27412 4924 27476 4928
rect 27412 4868 27416 4924
rect 27416 4868 27472 4924
rect 27472 4868 27476 4924
rect 27412 4864 27476 4868
rect 27492 4924 27556 4928
rect 27492 4868 27496 4924
rect 27496 4868 27552 4924
rect 27552 4868 27556 4924
rect 27492 4864 27556 4868
rect 1752 4380 1816 4384
rect 1752 4324 1756 4380
rect 1756 4324 1812 4380
rect 1812 4324 1816 4380
rect 1752 4320 1816 4324
rect 1832 4380 1896 4384
rect 1832 4324 1836 4380
rect 1836 4324 1892 4380
rect 1892 4324 1896 4380
rect 1832 4320 1896 4324
rect 1912 4380 1976 4384
rect 1912 4324 1916 4380
rect 1916 4324 1972 4380
rect 1972 4324 1976 4380
rect 1912 4320 1976 4324
rect 1992 4380 2056 4384
rect 1992 4324 1996 4380
rect 1996 4324 2052 4380
rect 2052 4324 2056 4380
rect 1992 4320 2056 4324
rect 4752 4380 4816 4384
rect 4752 4324 4756 4380
rect 4756 4324 4812 4380
rect 4812 4324 4816 4380
rect 4752 4320 4816 4324
rect 4832 4380 4896 4384
rect 4832 4324 4836 4380
rect 4836 4324 4892 4380
rect 4892 4324 4896 4380
rect 4832 4320 4896 4324
rect 4912 4380 4976 4384
rect 4912 4324 4916 4380
rect 4916 4324 4972 4380
rect 4972 4324 4976 4380
rect 4912 4320 4976 4324
rect 4992 4380 5056 4384
rect 4992 4324 4996 4380
rect 4996 4324 5052 4380
rect 5052 4324 5056 4380
rect 4992 4320 5056 4324
rect 7752 4380 7816 4384
rect 7752 4324 7756 4380
rect 7756 4324 7812 4380
rect 7812 4324 7816 4380
rect 7752 4320 7816 4324
rect 7832 4380 7896 4384
rect 7832 4324 7836 4380
rect 7836 4324 7892 4380
rect 7892 4324 7896 4380
rect 7832 4320 7896 4324
rect 7912 4380 7976 4384
rect 7912 4324 7916 4380
rect 7916 4324 7972 4380
rect 7972 4324 7976 4380
rect 7912 4320 7976 4324
rect 7992 4380 8056 4384
rect 7992 4324 7996 4380
rect 7996 4324 8052 4380
rect 8052 4324 8056 4380
rect 7992 4320 8056 4324
rect 10752 4380 10816 4384
rect 10752 4324 10756 4380
rect 10756 4324 10812 4380
rect 10812 4324 10816 4380
rect 10752 4320 10816 4324
rect 10832 4380 10896 4384
rect 10832 4324 10836 4380
rect 10836 4324 10892 4380
rect 10892 4324 10896 4380
rect 10832 4320 10896 4324
rect 10912 4380 10976 4384
rect 10912 4324 10916 4380
rect 10916 4324 10972 4380
rect 10972 4324 10976 4380
rect 10912 4320 10976 4324
rect 10992 4380 11056 4384
rect 10992 4324 10996 4380
rect 10996 4324 11052 4380
rect 11052 4324 11056 4380
rect 10992 4320 11056 4324
rect 13752 4380 13816 4384
rect 13752 4324 13756 4380
rect 13756 4324 13812 4380
rect 13812 4324 13816 4380
rect 13752 4320 13816 4324
rect 13832 4380 13896 4384
rect 13832 4324 13836 4380
rect 13836 4324 13892 4380
rect 13892 4324 13896 4380
rect 13832 4320 13896 4324
rect 13912 4380 13976 4384
rect 13912 4324 13916 4380
rect 13916 4324 13972 4380
rect 13972 4324 13976 4380
rect 13912 4320 13976 4324
rect 13992 4380 14056 4384
rect 13992 4324 13996 4380
rect 13996 4324 14052 4380
rect 14052 4324 14056 4380
rect 13992 4320 14056 4324
rect 16752 4380 16816 4384
rect 16752 4324 16756 4380
rect 16756 4324 16812 4380
rect 16812 4324 16816 4380
rect 16752 4320 16816 4324
rect 16832 4380 16896 4384
rect 16832 4324 16836 4380
rect 16836 4324 16892 4380
rect 16892 4324 16896 4380
rect 16832 4320 16896 4324
rect 16912 4380 16976 4384
rect 16912 4324 16916 4380
rect 16916 4324 16972 4380
rect 16972 4324 16976 4380
rect 16912 4320 16976 4324
rect 16992 4380 17056 4384
rect 16992 4324 16996 4380
rect 16996 4324 17052 4380
rect 17052 4324 17056 4380
rect 16992 4320 17056 4324
rect 19752 4380 19816 4384
rect 19752 4324 19756 4380
rect 19756 4324 19812 4380
rect 19812 4324 19816 4380
rect 19752 4320 19816 4324
rect 19832 4380 19896 4384
rect 19832 4324 19836 4380
rect 19836 4324 19892 4380
rect 19892 4324 19896 4380
rect 19832 4320 19896 4324
rect 19912 4380 19976 4384
rect 19912 4324 19916 4380
rect 19916 4324 19972 4380
rect 19972 4324 19976 4380
rect 19912 4320 19976 4324
rect 19992 4380 20056 4384
rect 19992 4324 19996 4380
rect 19996 4324 20052 4380
rect 20052 4324 20056 4380
rect 19992 4320 20056 4324
rect 22752 4380 22816 4384
rect 22752 4324 22756 4380
rect 22756 4324 22812 4380
rect 22812 4324 22816 4380
rect 22752 4320 22816 4324
rect 22832 4380 22896 4384
rect 22832 4324 22836 4380
rect 22836 4324 22892 4380
rect 22892 4324 22896 4380
rect 22832 4320 22896 4324
rect 22912 4380 22976 4384
rect 22912 4324 22916 4380
rect 22916 4324 22972 4380
rect 22972 4324 22976 4380
rect 22912 4320 22976 4324
rect 22992 4380 23056 4384
rect 22992 4324 22996 4380
rect 22996 4324 23052 4380
rect 23052 4324 23056 4380
rect 22992 4320 23056 4324
rect 25752 4380 25816 4384
rect 25752 4324 25756 4380
rect 25756 4324 25812 4380
rect 25812 4324 25816 4380
rect 25752 4320 25816 4324
rect 25832 4380 25896 4384
rect 25832 4324 25836 4380
rect 25836 4324 25892 4380
rect 25892 4324 25896 4380
rect 25832 4320 25896 4324
rect 25912 4380 25976 4384
rect 25912 4324 25916 4380
rect 25916 4324 25972 4380
rect 25972 4324 25976 4380
rect 25912 4320 25976 4324
rect 25992 4380 26056 4384
rect 25992 4324 25996 4380
rect 25996 4324 26052 4380
rect 26052 4324 26056 4380
rect 25992 4320 26056 4324
rect 3252 3836 3316 3840
rect 3252 3780 3256 3836
rect 3256 3780 3312 3836
rect 3312 3780 3316 3836
rect 3252 3776 3316 3780
rect 3332 3836 3396 3840
rect 3332 3780 3336 3836
rect 3336 3780 3392 3836
rect 3392 3780 3396 3836
rect 3332 3776 3396 3780
rect 3412 3836 3476 3840
rect 3412 3780 3416 3836
rect 3416 3780 3472 3836
rect 3472 3780 3476 3836
rect 3412 3776 3476 3780
rect 3492 3836 3556 3840
rect 3492 3780 3496 3836
rect 3496 3780 3552 3836
rect 3552 3780 3556 3836
rect 3492 3776 3556 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 6412 3836 6476 3840
rect 6412 3780 6416 3836
rect 6416 3780 6472 3836
rect 6472 3780 6476 3836
rect 6412 3776 6476 3780
rect 6492 3836 6556 3840
rect 6492 3780 6496 3836
rect 6496 3780 6552 3836
rect 6552 3780 6556 3836
rect 6492 3776 6556 3780
rect 9252 3836 9316 3840
rect 9252 3780 9256 3836
rect 9256 3780 9312 3836
rect 9312 3780 9316 3836
rect 9252 3776 9316 3780
rect 9332 3836 9396 3840
rect 9332 3780 9336 3836
rect 9336 3780 9392 3836
rect 9392 3780 9396 3836
rect 9332 3776 9396 3780
rect 9412 3836 9476 3840
rect 9412 3780 9416 3836
rect 9416 3780 9472 3836
rect 9472 3780 9476 3836
rect 9412 3776 9476 3780
rect 9492 3836 9556 3840
rect 9492 3780 9496 3836
rect 9496 3780 9552 3836
rect 9552 3780 9556 3836
rect 9492 3776 9556 3780
rect 12252 3836 12316 3840
rect 12252 3780 12256 3836
rect 12256 3780 12312 3836
rect 12312 3780 12316 3836
rect 12252 3776 12316 3780
rect 12332 3836 12396 3840
rect 12332 3780 12336 3836
rect 12336 3780 12392 3836
rect 12392 3780 12396 3836
rect 12332 3776 12396 3780
rect 12412 3836 12476 3840
rect 12412 3780 12416 3836
rect 12416 3780 12472 3836
rect 12472 3780 12476 3836
rect 12412 3776 12476 3780
rect 12492 3836 12556 3840
rect 12492 3780 12496 3836
rect 12496 3780 12552 3836
rect 12552 3780 12556 3836
rect 12492 3776 12556 3780
rect 15252 3836 15316 3840
rect 15252 3780 15256 3836
rect 15256 3780 15312 3836
rect 15312 3780 15316 3836
rect 15252 3776 15316 3780
rect 15332 3836 15396 3840
rect 15332 3780 15336 3836
rect 15336 3780 15392 3836
rect 15392 3780 15396 3836
rect 15332 3776 15396 3780
rect 15412 3836 15476 3840
rect 15412 3780 15416 3836
rect 15416 3780 15472 3836
rect 15472 3780 15476 3836
rect 15412 3776 15476 3780
rect 15492 3836 15556 3840
rect 15492 3780 15496 3836
rect 15496 3780 15552 3836
rect 15552 3780 15556 3836
rect 15492 3776 15556 3780
rect 18252 3836 18316 3840
rect 18252 3780 18256 3836
rect 18256 3780 18312 3836
rect 18312 3780 18316 3836
rect 18252 3776 18316 3780
rect 18332 3836 18396 3840
rect 18332 3780 18336 3836
rect 18336 3780 18392 3836
rect 18392 3780 18396 3836
rect 18332 3776 18396 3780
rect 18412 3836 18476 3840
rect 18412 3780 18416 3836
rect 18416 3780 18472 3836
rect 18472 3780 18476 3836
rect 18412 3776 18476 3780
rect 18492 3836 18556 3840
rect 18492 3780 18496 3836
rect 18496 3780 18552 3836
rect 18552 3780 18556 3836
rect 18492 3776 18556 3780
rect 21252 3836 21316 3840
rect 21252 3780 21256 3836
rect 21256 3780 21312 3836
rect 21312 3780 21316 3836
rect 21252 3776 21316 3780
rect 21332 3836 21396 3840
rect 21332 3780 21336 3836
rect 21336 3780 21392 3836
rect 21392 3780 21396 3836
rect 21332 3776 21396 3780
rect 21412 3836 21476 3840
rect 21412 3780 21416 3836
rect 21416 3780 21472 3836
rect 21472 3780 21476 3836
rect 21412 3776 21476 3780
rect 21492 3836 21556 3840
rect 21492 3780 21496 3836
rect 21496 3780 21552 3836
rect 21552 3780 21556 3836
rect 21492 3776 21556 3780
rect 24252 3836 24316 3840
rect 24252 3780 24256 3836
rect 24256 3780 24312 3836
rect 24312 3780 24316 3836
rect 24252 3776 24316 3780
rect 24332 3836 24396 3840
rect 24332 3780 24336 3836
rect 24336 3780 24392 3836
rect 24392 3780 24396 3836
rect 24332 3776 24396 3780
rect 24412 3836 24476 3840
rect 24412 3780 24416 3836
rect 24416 3780 24472 3836
rect 24472 3780 24476 3836
rect 24412 3776 24476 3780
rect 24492 3836 24556 3840
rect 24492 3780 24496 3836
rect 24496 3780 24552 3836
rect 24552 3780 24556 3836
rect 24492 3776 24556 3780
rect 27252 3836 27316 3840
rect 27252 3780 27256 3836
rect 27256 3780 27312 3836
rect 27312 3780 27316 3836
rect 27252 3776 27316 3780
rect 27332 3836 27396 3840
rect 27332 3780 27336 3836
rect 27336 3780 27392 3836
rect 27392 3780 27396 3836
rect 27332 3776 27396 3780
rect 27412 3836 27476 3840
rect 27412 3780 27416 3836
rect 27416 3780 27472 3836
rect 27472 3780 27476 3836
rect 27412 3776 27476 3780
rect 27492 3836 27556 3840
rect 27492 3780 27496 3836
rect 27496 3780 27552 3836
rect 27552 3780 27556 3836
rect 27492 3776 27556 3780
rect 1752 3292 1816 3296
rect 1752 3236 1756 3292
rect 1756 3236 1812 3292
rect 1812 3236 1816 3292
rect 1752 3232 1816 3236
rect 1832 3292 1896 3296
rect 1832 3236 1836 3292
rect 1836 3236 1892 3292
rect 1892 3236 1896 3292
rect 1832 3232 1896 3236
rect 1912 3292 1976 3296
rect 1912 3236 1916 3292
rect 1916 3236 1972 3292
rect 1972 3236 1976 3292
rect 1912 3232 1976 3236
rect 1992 3292 2056 3296
rect 1992 3236 1996 3292
rect 1996 3236 2052 3292
rect 2052 3236 2056 3292
rect 1992 3232 2056 3236
rect 4752 3292 4816 3296
rect 4752 3236 4756 3292
rect 4756 3236 4812 3292
rect 4812 3236 4816 3292
rect 4752 3232 4816 3236
rect 4832 3292 4896 3296
rect 4832 3236 4836 3292
rect 4836 3236 4892 3292
rect 4892 3236 4896 3292
rect 4832 3232 4896 3236
rect 4912 3292 4976 3296
rect 4912 3236 4916 3292
rect 4916 3236 4972 3292
rect 4972 3236 4976 3292
rect 4912 3232 4976 3236
rect 4992 3292 5056 3296
rect 4992 3236 4996 3292
rect 4996 3236 5052 3292
rect 5052 3236 5056 3292
rect 4992 3232 5056 3236
rect 7752 3292 7816 3296
rect 7752 3236 7756 3292
rect 7756 3236 7812 3292
rect 7812 3236 7816 3292
rect 7752 3232 7816 3236
rect 7832 3292 7896 3296
rect 7832 3236 7836 3292
rect 7836 3236 7892 3292
rect 7892 3236 7896 3292
rect 7832 3232 7896 3236
rect 7912 3292 7976 3296
rect 7912 3236 7916 3292
rect 7916 3236 7972 3292
rect 7972 3236 7976 3292
rect 7912 3232 7976 3236
rect 7992 3292 8056 3296
rect 7992 3236 7996 3292
rect 7996 3236 8052 3292
rect 8052 3236 8056 3292
rect 7992 3232 8056 3236
rect 10752 3292 10816 3296
rect 10752 3236 10756 3292
rect 10756 3236 10812 3292
rect 10812 3236 10816 3292
rect 10752 3232 10816 3236
rect 10832 3292 10896 3296
rect 10832 3236 10836 3292
rect 10836 3236 10892 3292
rect 10892 3236 10896 3292
rect 10832 3232 10896 3236
rect 10912 3292 10976 3296
rect 10912 3236 10916 3292
rect 10916 3236 10972 3292
rect 10972 3236 10976 3292
rect 10912 3232 10976 3236
rect 10992 3292 11056 3296
rect 10992 3236 10996 3292
rect 10996 3236 11052 3292
rect 11052 3236 11056 3292
rect 10992 3232 11056 3236
rect 13752 3292 13816 3296
rect 13752 3236 13756 3292
rect 13756 3236 13812 3292
rect 13812 3236 13816 3292
rect 13752 3232 13816 3236
rect 13832 3292 13896 3296
rect 13832 3236 13836 3292
rect 13836 3236 13892 3292
rect 13892 3236 13896 3292
rect 13832 3232 13896 3236
rect 13912 3292 13976 3296
rect 13912 3236 13916 3292
rect 13916 3236 13972 3292
rect 13972 3236 13976 3292
rect 13912 3232 13976 3236
rect 13992 3292 14056 3296
rect 13992 3236 13996 3292
rect 13996 3236 14052 3292
rect 14052 3236 14056 3292
rect 13992 3232 14056 3236
rect 16752 3292 16816 3296
rect 16752 3236 16756 3292
rect 16756 3236 16812 3292
rect 16812 3236 16816 3292
rect 16752 3232 16816 3236
rect 16832 3292 16896 3296
rect 16832 3236 16836 3292
rect 16836 3236 16892 3292
rect 16892 3236 16896 3292
rect 16832 3232 16896 3236
rect 16912 3292 16976 3296
rect 16912 3236 16916 3292
rect 16916 3236 16972 3292
rect 16972 3236 16976 3292
rect 16912 3232 16976 3236
rect 16992 3292 17056 3296
rect 16992 3236 16996 3292
rect 16996 3236 17052 3292
rect 17052 3236 17056 3292
rect 16992 3232 17056 3236
rect 19752 3292 19816 3296
rect 19752 3236 19756 3292
rect 19756 3236 19812 3292
rect 19812 3236 19816 3292
rect 19752 3232 19816 3236
rect 19832 3292 19896 3296
rect 19832 3236 19836 3292
rect 19836 3236 19892 3292
rect 19892 3236 19896 3292
rect 19832 3232 19896 3236
rect 19912 3292 19976 3296
rect 19912 3236 19916 3292
rect 19916 3236 19972 3292
rect 19972 3236 19976 3292
rect 19912 3232 19976 3236
rect 19992 3292 20056 3296
rect 19992 3236 19996 3292
rect 19996 3236 20052 3292
rect 20052 3236 20056 3292
rect 19992 3232 20056 3236
rect 22752 3292 22816 3296
rect 22752 3236 22756 3292
rect 22756 3236 22812 3292
rect 22812 3236 22816 3292
rect 22752 3232 22816 3236
rect 22832 3292 22896 3296
rect 22832 3236 22836 3292
rect 22836 3236 22892 3292
rect 22892 3236 22896 3292
rect 22832 3232 22896 3236
rect 22912 3292 22976 3296
rect 22912 3236 22916 3292
rect 22916 3236 22972 3292
rect 22972 3236 22976 3292
rect 22912 3232 22976 3236
rect 22992 3292 23056 3296
rect 22992 3236 22996 3292
rect 22996 3236 23052 3292
rect 23052 3236 23056 3292
rect 22992 3232 23056 3236
rect 25752 3292 25816 3296
rect 25752 3236 25756 3292
rect 25756 3236 25812 3292
rect 25812 3236 25816 3292
rect 25752 3232 25816 3236
rect 25832 3292 25896 3296
rect 25832 3236 25836 3292
rect 25836 3236 25892 3292
rect 25892 3236 25896 3292
rect 25832 3232 25896 3236
rect 25912 3292 25976 3296
rect 25912 3236 25916 3292
rect 25916 3236 25972 3292
rect 25972 3236 25976 3292
rect 25912 3232 25976 3236
rect 25992 3292 26056 3296
rect 25992 3236 25996 3292
rect 25996 3236 26052 3292
rect 26052 3236 26056 3292
rect 25992 3232 26056 3236
rect 3252 2748 3316 2752
rect 3252 2692 3256 2748
rect 3256 2692 3312 2748
rect 3312 2692 3316 2748
rect 3252 2688 3316 2692
rect 3332 2748 3396 2752
rect 3332 2692 3336 2748
rect 3336 2692 3392 2748
rect 3392 2692 3396 2748
rect 3332 2688 3396 2692
rect 3412 2748 3476 2752
rect 3412 2692 3416 2748
rect 3416 2692 3472 2748
rect 3472 2692 3476 2748
rect 3412 2688 3476 2692
rect 3492 2748 3556 2752
rect 3492 2692 3496 2748
rect 3496 2692 3552 2748
rect 3552 2692 3556 2748
rect 3492 2688 3556 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 6412 2748 6476 2752
rect 6412 2692 6416 2748
rect 6416 2692 6472 2748
rect 6472 2692 6476 2748
rect 6412 2688 6476 2692
rect 6492 2748 6556 2752
rect 6492 2692 6496 2748
rect 6496 2692 6552 2748
rect 6552 2692 6556 2748
rect 6492 2688 6556 2692
rect 9252 2748 9316 2752
rect 9252 2692 9256 2748
rect 9256 2692 9312 2748
rect 9312 2692 9316 2748
rect 9252 2688 9316 2692
rect 9332 2748 9396 2752
rect 9332 2692 9336 2748
rect 9336 2692 9392 2748
rect 9392 2692 9396 2748
rect 9332 2688 9396 2692
rect 9412 2748 9476 2752
rect 9412 2692 9416 2748
rect 9416 2692 9472 2748
rect 9472 2692 9476 2748
rect 9412 2688 9476 2692
rect 9492 2748 9556 2752
rect 9492 2692 9496 2748
rect 9496 2692 9552 2748
rect 9552 2692 9556 2748
rect 9492 2688 9556 2692
rect 12252 2748 12316 2752
rect 12252 2692 12256 2748
rect 12256 2692 12312 2748
rect 12312 2692 12316 2748
rect 12252 2688 12316 2692
rect 12332 2748 12396 2752
rect 12332 2692 12336 2748
rect 12336 2692 12392 2748
rect 12392 2692 12396 2748
rect 12332 2688 12396 2692
rect 12412 2748 12476 2752
rect 12412 2692 12416 2748
rect 12416 2692 12472 2748
rect 12472 2692 12476 2748
rect 12412 2688 12476 2692
rect 12492 2748 12556 2752
rect 12492 2692 12496 2748
rect 12496 2692 12552 2748
rect 12552 2692 12556 2748
rect 12492 2688 12556 2692
rect 15252 2748 15316 2752
rect 15252 2692 15256 2748
rect 15256 2692 15312 2748
rect 15312 2692 15316 2748
rect 15252 2688 15316 2692
rect 15332 2748 15396 2752
rect 15332 2692 15336 2748
rect 15336 2692 15392 2748
rect 15392 2692 15396 2748
rect 15332 2688 15396 2692
rect 15412 2748 15476 2752
rect 15412 2692 15416 2748
rect 15416 2692 15472 2748
rect 15472 2692 15476 2748
rect 15412 2688 15476 2692
rect 15492 2748 15556 2752
rect 15492 2692 15496 2748
rect 15496 2692 15552 2748
rect 15552 2692 15556 2748
rect 15492 2688 15556 2692
rect 18252 2748 18316 2752
rect 18252 2692 18256 2748
rect 18256 2692 18312 2748
rect 18312 2692 18316 2748
rect 18252 2688 18316 2692
rect 18332 2748 18396 2752
rect 18332 2692 18336 2748
rect 18336 2692 18392 2748
rect 18392 2692 18396 2748
rect 18332 2688 18396 2692
rect 18412 2748 18476 2752
rect 18412 2692 18416 2748
rect 18416 2692 18472 2748
rect 18472 2692 18476 2748
rect 18412 2688 18476 2692
rect 18492 2748 18556 2752
rect 18492 2692 18496 2748
rect 18496 2692 18552 2748
rect 18552 2692 18556 2748
rect 18492 2688 18556 2692
rect 21252 2748 21316 2752
rect 21252 2692 21256 2748
rect 21256 2692 21312 2748
rect 21312 2692 21316 2748
rect 21252 2688 21316 2692
rect 21332 2748 21396 2752
rect 21332 2692 21336 2748
rect 21336 2692 21392 2748
rect 21392 2692 21396 2748
rect 21332 2688 21396 2692
rect 21412 2748 21476 2752
rect 21412 2692 21416 2748
rect 21416 2692 21472 2748
rect 21472 2692 21476 2748
rect 21412 2688 21476 2692
rect 21492 2748 21556 2752
rect 21492 2692 21496 2748
rect 21496 2692 21552 2748
rect 21552 2692 21556 2748
rect 21492 2688 21556 2692
rect 24252 2748 24316 2752
rect 24252 2692 24256 2748
rect 24256 2692 24312 2748
rect 24312 2692 24316 2748
rect 24252 2688 24316 2692
rect 24332 2748 24396 2752
rect 24332 2692 24336 2748
rect 24336 2692 24392 2748
rect 24392 2692 24396 2748
rect 24332 2688 24396 2692
rect 24412 2748 24476 2752
rect 24412 2692 24416 2748
rect 24416 2692 24472 2748
rect 24472 2692 24476 2748
rect 24412 2688 24476 2692
rect 24492 2748 24556 2752
rect 24492 2692 24496 2748
rect 24496 2692 24552 2748
rect 24552 2692 24556 2748
rect 24492 2688 24556 2692
rect 27252 2748 27316 2752
rect 27252 2692 27256 2748
rect 27256 2692 27312 2748
rect 27312 2692 27316 2748
rect 27252 2688 27316 2692
rect 27332 2748 27396 2752
rect 27332 2692 27336 2748
rect 27336 2692 27392 2748
rect 27392 2692 27396 2748
rect 27332 2688 27396 2692
rect 27412 2748 27476 2752
rect 27412 2692 27416 2748
rect 27416 2692 27472 2748
rect 27472 2692 27476 2748
rect 27412 2688 27476 2692
rect 27492 2748 27556 2752
rect 27492 2692 27496 2748
rect 27496 2692 27552 2748
rect 27552 2692 27556 2748
rect 27492 2688 27556 2692
rect 1752 2204 1816 2208
rect 1752 2148 1756 2204
rect 1756 2148 1812 2204
rect 1812 2148 1816 2204
rect 1752 2144 1816 2148
rect 1832 2204 1896 2208
rect 1832 2148 1836 2204
rect 1836 2148 1892 2204
rect 1892 2148 1896 2204
rect 1832 2144 1896 2148
rect 1912 2204 1976 2208
rect 1912 2148 1916 2204
rect 1916 2148 1972 2204
rect 1972 2148 1976 2204
rect 1912 2144 1976 2148
rect 1992 2204 2056 2208
rect 1992 2148 1996 2204
rect 1996 2148 2052 2204
rect 2052 2148 2056 2204
rect 1992 2144 2056 2148
rect 4752 2204 4816 2208
rect 4752 2148 4756 2204
rect 4756 2148 4812 2204
rect 4812 2148 4816 2204
rect 4752 2144 4816 2148
rect 4832 2204 4896 2208
rect 4832 2148 4836 2204
rect 4836 2148 4892 2204
rect 4892 2148 4896 2204
rect 4832 2144 4896 2148
rect 4912 2204 4976 2208
rect 4912 2148 4916 2204
rect 4916 2148 4972 2204
rect 4972 2148 4976 2204
rect 4912 2144 4976 2148
rect 4992 2204 5056 2208
rect 4992 2148 4996 2204
rect 4996 2148 5052 2204
rect 5052 2148 5056 2204
rect 4992 2144 5056 2148
rect 7752 2204 7816 2208
rect 7752 2148 7756 2204
rect 7756 2148 7812 2204
rect 7812 2148 7816 2204
rect 7752 2144 7816 2148
rect 7832 2204 7896 2208
rect 7832 2148 7836 2204
rect 7836 2148 7892 2204
rect 7892 2148 7896 2204
rect 7832 2144 7896 2148
rect 7912 2204 7976 2208
rect 7912 2148 7916 2204
rect 7916 2148 7972 2204
rect 7972 2148 7976 2204
rect 7912 2144 7976 2148
rect 7992 2204 8056 2208
rect 7992 2148 7996 2204
rect 7996 2148 8052 2204
rect 8052 2148 8056 2204
rect 7992 2144 8056 2148
rect 10752 2204 10816 2208
rect 10752 2148 10756 2204
rect 10756 2148 10812 2204
rect 10812 2148 10816 2204
rect 10752 2144 10816 2148
rect 10832 2204 10896 2208
rect 10832 2148 10836 2204
rect 10836 2148 10892 2204
rect 10892 2148 10896 2204
rect 10832 2144 10896 2148
rect 10912 2204 10976 2208
rect 10912 2148 10916 2204
rect 10916 2148 10972 2204
rect 10972 2148 10976 2204
rect 10912 2144 10976 2148
rect 10992 2204 11056 2208
rect 10992 2148 10996 2204
rect 10996 2148 11052 2204
rect 11052 2148 11056 2204
rect 10992 2144 11056 2148
rect 13752 2204 13816 2208
rect 13752 2148 13756 2204
rect 13756 2148 13812 2204
rect 13812 2148 13816 2204
rect 13752 2144 13816 2148
rect 13832 2204 13896 2208
rect 13832 2148 13836 2204
rect 13836 2148 13892 2204
rect 13892 2148 13896 2204
rect 13832 2144 13896 2148
rect 13912 2204 13976 2208
rect 13912 2148 13916 2204
rect 13916 2148 13972 2204
rect 13972 2148 13976 2204
rect 13912 2144 13976 2148
rect 13992 2204 14056 2208
rect 13992 2148 13996 2204
rect 13996 2148 14052 2204
rect 14052 2148 14056 2204
rect 13992 2144 14056 2148
rect 16752 2204 16816 2208
rect 16752 2148 16756 2204
rect 16756 2148 16812 2204
rect 16812 2148 16816 2204
rect 16752 2144 16816 2148
rect 16832 2204 16896 2208
rect 16832 2148 16836 2204
rect 16836 2148 16892 2204
rect 16892 2148 16896 2204
rect 16832 2144 16896 2148
rect 16912 2204 16976 2208
rect 16912 2148 16916 2204
rect 16916 2148 16972 2204
rect 16972 2148 16976 2204
rect 16912 2144 16976 2148
rect 16992 2204 17056 2208
rect 16992 2148 16996 2204
rect 16996 2148 17052 2204
rect 17052 2148 17056 2204
rect 16992 2144 17056 2148
rect 19752 2204 19816 2208
rect 19752 2148 19756 2204
rect 19756 2148 19812 2204
rect 19812 2148 19816 2204
rect 19752 2144 19816 2148
rect 19832 2204 19896 2208
rect 19832 2148 19836 2204
rect 19836 2148 19892 2204
rect 19892 2148 19896 2204
rect 19832 2144 19896 2148
rect 19912 2204 19976 2208
rect 19912 2148 19916 2204
rect 19916 2148 19972 2204
rect 19972 2148 19976 2204
rect 19912 2144 19976 2148
rect 19992 2204 20056 2208
rect 19992 2148 19996 2204
rect 19996 2148 20052 2204
rect 20052 2148 20056 2204
rect 19992 2144 20056 2148
rect 22752 2204 22816 2208
rect 22752 2148 22756 2204
rect 22756 2148 22812 2204
rect 22812 2148 22816 2204
rect 22752 2144 22816 2148
rect 22832 2204 22896 2208
rect 22832 2148 22836 2204
rect 22836 2148 22892 2204
rect 22892 2148 22896 2204
rect 22832 2144 22896 2148
rect 22912 2204 22976 2208
rect 22912 2148 22916 2204
rect 22916 2148 22972 2204
rect 22972 2148 22976 2204
rect 22912 2144 22976 2148
rect 22992 2204 23056 2208
rect 22992 2148 22996 2204
rect 22996 2148 23052 2204
rect 23052 2148 23056 2204
rect 22992 2144 23056 2148
rect 25752 2204 25816 2208
rect 25752 2148 25756 2204
rect 25756 2148 25812 2204
rect 25812 2148 25816 2204
rect 25752 2144 25816 2148
rect 25832 2204 25896 2208
rect 25832 2148 25836 2204
rect 25836 2148 25892 2204
rect 25892 2148 25896 2204
rect 25832 2144 25896 2148
rect 25912 2204 25976 2208
rect 25912 2148 25916 2204
rect 25916 2148 25972 2204
rect 25972 2148 25976 2204
rect 25912 2144 25976 2148
rect 25992 2204 26056 2208
rect 25992 2148 25996 2204
rect 25996 2148 26052 2204
rect 26052 2148 26056 2204
rect 25992 2144 26056 2148
<< metal4 >>
rect 1744 29408 2064 29424
rect 1744 29344 1752 29408
rect 1816 29344 1832 29408
rect 1896 29344 1912 29408
rect 1976 29344 1992 29408
rect 2056 29344 2064 29408
rect 1744 28320 2064 29344
rect 1744 28256 1752 28320
rect 1816 28256 1832 28320
rect 1896 28256 1912 28320
rect 1976 28256 1992 28320
rect 2056 28256 2064 28320
rect 1744 27232 2064 28256
rect 1744 27168 1752 27232
rect 1816 27168 1832 27232
rect 1896 27168 1912 27232
rect 1976 27168 1992 27232
rect 2056 27168 2064 27232
rect 1744 27046 2064 27168
rect 1744 26810 1786 27046
rect 2022 26810 2064 27046
rect 1744 26144 2064 26810
rect 1744 26080 1752 26144
rect 1816 26080 1832 26144
rect 1896 26080 1912 26144
rect 1976 26080 1992 26144
rect 2056 26080 2064 26144
rect 1744 25056 2064 26080
rect 1744 24992 1752 25056
rect 1816 24992 1832 25056
rect 1896 24992 1912 25056
rect 1976 24992 1992 25056
rect 2056 24992 2064 25056
rect 1744 24046 2064 24992
rect 1744 23968 1786 24046
rect 2022 23968 2064 24046
rect 1744 23904 1752 23968
rect 2056 23904 2064 23968
rect 1744 23810 1786 23904
rect 2022 23810 2064 23904
rect 1744 22880 2064 23810
rect 1744 22816 1752 22880
rect 1816 22816 1832 22880
rect 1896 22816 1912 22880
rect 1976 22816 1992 22880
rect 2056 22816 2064 22880
rect 1744 21792 2064 22816
rect 1744 21728 1752 21792
rect 1816 21728 1832 21792
rect 1896 21728 1912 21792
rect 1976 21728 1992 21792
rect 2056 21728 2064 21792
rect 1744 21046 2064 21728
rect 1744 20810 1786 21046
rect 2022 20810 2064 21046
rect 1744 20704 2064 20810
rect 1744 20640 1752 20704
rect 1816 20640 1832 20704
rect 1896 20640 1912 20704
rect 1976 20640 1992 20704
rect 2056 20640 2064 20704
rect 1744 19616 2064 20640
rect 1744 19552 1752 19616
rect 1816 19552 1832 19616
rect 1896 19552 1912 19616
rect 1976 19552 1992 19616
rect 2056 19552 2064 19616
rect 1744 18528 2064 19552
rect 1744 18464 1752 18528
rect 1816 18464 1832 18528
rect 1896 18464 1912 18528
rect 1976 18464 1992 18528
rect 2056 18464 2064 18528
rect 1744 18046 2064 18464
rect 1744 17810 1786 18046
rect 2022 17810 2064 18046
rect 1744 17440 2064 17810
rect 1744 17376 1752 17440
rect 1816 17376 1832 17440
rect 1896 17376 1912 17440
rect 1976 17376 1992 17440
rect 2056 17376 2064 17440
rect 1744 16352 2064 17376
rect 1744 16288 1752 16352
rect 1816 16288 1832 16352
rect 1896 16288 1912 16352
rect 1976 16288 1992 16352
rect 2056 16288 2064 16352
rect 1744 15264 2064 16288
rect 1744 15200 1752 15264
rect 1816 15200 1832 15264
rect 1896 15200 1912 15264
rect 1976 15200 1992 15264
rect 2056 15200 2064 15264
rect 1744 15046 2064 15200
rect 1744 14810 1786 15046
rect 2022 14810 2064 15046
rect 1744 14176 2064 14810
rect 1744 14112 1752 14176
rect 1816 14112 1832 14176
rect 1896 14112 1912 14176
rect 1976 14112 1992 14176
rect 2056 14112 2064 14176
rect 1744 13088 2064 14112
rect 1744 13024 1752 13088
rect 1816 13024 1832 13088
rect 1896 13024 1912 13088
rect 1976 13024 1992 13088
rect 2056 13024 2064 13088
rect 1744 12046 2064 13024
rect 1744 12000 1786 12046
rect 2022 12000 2064 12046
rect 1744 11936 1752 12000
rect 2056 11936 2064 12000
rect 1744 11810 1786 11936
rect 2022 11810 2064 11936
rect 1744 10912 2064 11810
rect 1744 10848 1752 10912
rect 1816 10848 1832 10912
rect 1896 10848 1912 10912
rect 1976 10848 1992 10912
rect 2056 10848 2064 10912
rect 1744 9824 2064 10848
rect 1744 9760 1752 9824
rect 1816 9760 1832 9824
rect 1896 9760 1912 9824
rect 1976 9760 1992 9824
rect 2056 9760 2064 9824
rect 1744 9046 2064 9760
rect 1744 8810 1786 9046
rect 2022 8810 2064 9046
rect 1744 8736 2064 8810
rect 1744 8672 1752 8736
rect 1816 8672 1832 8736
rect 1896 8672 1912 8736
rect 1976 8672 1992 8736
rect 2056 8672 2064 8736
rect 1744 7648 2064 8672
rect 1744 7584 1752 7648
rect 1816 7584 1832 7648
rect 1896 7584 1912 7648
rect 1976 7584 1992 7648
rect 2056 7584 2064 7648
rect 1744 6560 2064 7584
rect 1744 6496 1752 6560
rect 1816 6496 1832 6560
rect 1896 6496 1912 6560
rect 1976 6496 1992 6560
rect 2056 6496 2064 6560
rect 1744 6046 2064 6496
rect 1744 5810 1786 6046
rect 2022 5810 2064 6046
rect 1744 5472 2064 5810
rect 1744 5408 1752 5472
rect 1816 5408 1832 5472
rect 1896 5408 1912 5472
rect 1976 5408 1992 5472
rect 2056 5408 2064 5472
rect 1744 4384 2064 5408
rect 1744 4320 1752 4384
rect 1816 4320 1832 4384
rect 1896 4320 1912 4384
rect 1976 4320 1992 4384
rect 2056 4320 2064 4384
rect 1744 3296 2064 4320
rect 1744 3232 1752 3296
rect 1816 3232 1832 3296
rect 1896 3232 1912 3296
rect 1976 3232 1992 3296
rect 2056 3232 2064 3296
rect 1744 3046 2064 3232
rect 1744 2810 1786 3046
rect 2022 2810 2064 3046
rect 1744 2208 2064 2810
rect 1744 2144 1752 2208
rect 1816 2144 1832 2208
rect 1896 2144 1912 2208
rect 1976 2144 1992 2208
rect 2056 2144 2064 2208
rect 1744 2128 2064 2144
rect 3244 28864 3564 29424
rect 3244 28800 3252 28864
rect 3316 28800 3332 28864
rect 3396 28800 3412 28864
rect 3476 28800 3492 28864
rect 3556 28800 3564 28864
rect 3244 28546 3564 28800
rect 3244 28310 3286 28546
rect 3522 28310 3564 28546
rect 3244 27776 3564 28310
rect 3244 27712 3252 27776
rect 3316 27712 3332 27776
rect 3396 27712 3412 27776
rect 3476 27712 3492 27776
rect 3556 27712 3564 27776
rect 3244 26688 3564 27712
rect 3244 26624 3252 26688
rect 3316 26624 3332 26688
rect 3396 26624 3412 26688
rect 3476 26624 3492 26688
rect 3556 26624 3564 26688
rect 3244 25600 3564 26624
rect 3244 25536 3252 25600
rect 3316 25546 3332 25600
rect 3396 25546 3412 25600
rect 3476 25546 3492 25600
rect 3556 25536 3564 25600
rect 3244 25310 3286 25536
rect 3522 25310 3564 25536
rect 3244 24512 3564 25310
rect 3244 24448 3252 24512
rect 3316 24448 3332 24512
rect 3396 24448 3412 24512
rect 3476 24448 3492 24512
rect 3556 24448 3564 24512
rect 3244 23424 3564 24448
rect 3244 23360 3252 23424
rect 3316 23360 3332 23424
rect 3396 23360 3412 23424
rect 3476 23360 3492 23424
rect 3556 23360 3564 23424
rect 3244 22546 3564 23360
rect 3244 22336 3286 22546
rect 3522 22336 3564 22546
rect 3244 22272 3252 22336
rect 3316 22272 3332 22310
rect 3396 22272 3412 22310
rect 3476 22272 3492 22310
rect 3556 22272 3564 22336
rect 3244 21248 3564 22272
rect 3244 21184 3252 21248
rect 3316 21184 3332 21248
rect 3396 21184 3412 21248
rect 3476 21184 3492 21248
rect 3556 21184 3564 21248
rect 3244 20160 3564 21184
rect 3244 20096 3252 20160
rect 3316 20096 3332 20160
rect 3396 20096 3412 20160
rect 3476 20096 3492 20160
rect 3556 20096 3564 20160
rect 3244 19546 3564 20096
rect 3244 19310 3286 19546
rect 3522 19310 3564 19546
rect 3244 19072 3564 19310
rect 3244 19008 3252 19072
rect 3316 19008 3332 19072
rect 3396 19008 3412 19072
rect 3476 19008 3492 19072
rect 3556 19008 3564 19072
rect 3244 17984 3564 19008
rect 3244 17920 3252 17984
rect 3316 17920 3332 17984
rect 3396 17920 3412 17984
rect 3476 17920 3492 17984
rect 3556 17920 3564 17984
rect 3244 16896 3564 17920
rect 3244 16832 3252 16896
rect 3316 16832 3332 16896
rect 3396 16832 3412 16896
rect 3476 16832 3492 16896
rect 3556 16832 3564 16896
rect 3244 16546 3564 16832
rect 3244 16310 3286 16546
rect 3522 16310 3564 16546
rect 3244 15808 3564 16310
rect 3244 15744 3252 15808
rect 3316 15744 3332 15808
rect 3396 15744 3412 15808
rect 3476 15744 3492 15808
rect 3556 15744 3564 15808
rect 3244 14720 3564 15744
rect 3244 14656 3252 14720
rect 3316 14656 3332 14720
rect 3396 14656 3412 14720
rect 3476 14656 3492 14720
rect 3556 14656 3564 14720
rect 3244 13632 3564 14656
rect 3244 13568 3252 13632
rect 3316 13568 3332 13632
rect 3396 13568 3412 13632
rect 3476 13568 3492 13632
rect 3556 13568 3564 13632
rect 3244 13546 3564 13568
rect 3244 13310 3286 13546
rect 3522 13310 3564 13546
rect 3244 12544 3564 13310
rect 3244 12480 3252 12544
rect 3316 12480 3332 12544
rect 3396 12480 3412 12544
rect 3476 12480 3492 12544
rect 3556 12480 3564 12544
rect 3244 11456 3564 12480
rect 3244 11392 3252 11456
rect 3316 11392 3332 11456
rect 3396 11392 3412 11456
rect 3476 11392 3492 11456
rect 3556 11392 3564 11456
rect 3244 10546 3564 11392
rect 3244 10368 3286 10546
rect 3522 10368 3564 10546
rect 3244 10304 3252 10368
rect 3316 10304 3332 10310
rect 3396 10304 3412 10310
rect 3476 10304 3492 10310
rect 3556 10304 3564 10368
rect 3244 9280 3564 10304
rect 3244 9216 3252 9280
rect 3316 9216 3332 9280
rect 3396 9216 3412 9280
rect 3476 9216 3492 9280
rect 3556 9216 3564 9280
rect 3244 8192 3564 9216
rect 3244 8128 3252 8192
rect 3316 8128 3332 8192
rect 3396 8128 3412 8192
rect 3476 8128 3492 8192
rect 3556 8128 3564 8192
rect 3244 7546 3564 8128
rect 3244 7310 3286 7546
rect 3522 7310 3564 7546
rect 3244 7104 3564 7310
rect 3244 7040 3252 7104
rect 3316 7040 3332 7104
rect 3396 7040 3412 7104
rect 3476 7040 3492 7104
rect 3556 7040 3564 7104
rect 3244 6016 3564 7040
rect 3244 5952 3252 6016
rect 3316 5952 3332 6016
rect 3396 5952 3412 6016
rect 3476 5952 3492 6016
rect 3556 5952 3564 6016
rect 3244 4928 3564 5952
rect 3244 4864 3252 4928
rect 3316 4864 3332 4928
rect 3396 4864 3412 4928
rect 3476 4864 3492 4928
rect 3556 4864 3564 4928
rect 3244 4546 3564 4864
rect 3244 4310 3286 4546
rect 3522 4310 3564 4546
rect 3244 3840 3564 4310
rect 3244 3776 3252 3840
rect 3316 3776 3332 3840
rect 3396 3776 3412 3840
rect 3476 3776 3492 3840
rect 3556 3776 3564 3840
rect 3244 2752 3564 3776
rect 3244 2688 3252 2752
rect 3316 2688 3332 2752
rect 3396 2688 3412 2752
rect 3476 2688 3492 2752
rect 3556 2688 3564 2752
rect 3244 2128 3564 2688
rect 4744 29408 5064 29424
rect 4744 29344 4752 29408
rect 4816 29344 4832 29408
rect 4896 29344 4912 29408
rect 4976 29344 4992 29408
rect 5056 29344 5064 29408
rect 4744 28320 5064 29344
rect 4744 28256 4752 28320
rect 4816 28256 4832 28320
rect 4896 28256 4912 28320
rect 4976 28256 4992 28320
rect 5056 28256 5064 28320
rect 4744 27232 5064 28256
rect 4744 27168 4752 27232
rect 4816 27168 4832 27232
rect 4896 27168 4912 27232
rect 4976 27168 4992 27232
rect 5056 27168 5064 27232
rect 4744 27046 5064 27168
rect 4744 26810 4786 27046
rect 5022 26810 5064 27046
rect 4744 26144 5064 26810
rect 4744 26080 4752 26144
rect 4816 26080 4832 26144
rect 4896 26080 4912 26144
rect 4976 26080 4992 26144
rect 5056 26080 5064 26144
rect 4744 25056 5064 26080
rect 4744 24992 4752 25056
rect 4816 24992 4832 25056
rect 4896 24992 4912 25056
rect 4976 24992 4992 25056
rect 5056 24992 5064 25056
rect 4744 24046 5064 24992
rect 4744 23968 4786 24046
rect 5022 23968 5064 24046
rect 4744 23904 4752 23968
rect 5056 23904 5064 23968
rect 4744 23810 4786 23904
rect 5022 23810 5064 23904
rect 4744 22880 5064 23810
rect 4744 22816 4752 22880
rect 4816 22816 4832 22880
rect 4896 22816 4912 22880
rect 4976 22816 4992 22880
rect 5056 22816 5064 22880
rect 4744 21792 5064 22816
rect 4744 21728 4752 21792
rect 4816 21728 4832 21792
rect 4896 21728 4912 21792
rect 4976 21728 4992 21792
rect 5056 21728 5064 21792
rect 4744 21046 5064 21728
rect 4744 20810 4786 21046
rect 5022 20810 5064 21046
rect 4744 20704 5064 20810
rect 4744 20640 4752 20704
rect 4816 20640 4832 20704
rect 4896 20640 4912 20704
rect 4976 20640 4992 20704
rect 5056 20640 5064 20704
rect 4744 19616 5064 20640
rect 4744 19552 4752 19616
rect 4816 19552 4832 19616
rect 4896 19552 4912 19616
rect 4976 19552 4992 19616
rect 5056 19552 5064 19616
rect 4744 18528 5064 19552
rect 4744 18464 4752 18528
rect 4816 18464 4832 18528
rect 4896 18464 4912 18528
rect 4976 18464 4992 18528
rect 5056 18464 5064 18528
rect 4744 18046 5064 18464
rect 4744 17810 4786 18046
rect 5022 17810 5064 18046
rect 4744 17440 5064 17810
rect 4744 17376 4752 17440
rect 4816 17376 4832 17440
rect 4896 17376 4912 17440
rect 4976 17376 4992 17440
rect 5056 17376 5064 17440
rect 4744 16352 5064 17376
rect 4744 16288 4752 16352
rect 4816 16288 4832 16352
rect 4896 16288 4912 16352
rect 4976 16288 4992 16352
rect 5056 16288 5064 16352
rect 4744 15264 5064 16288
rect 4744 15200 4752 15264
rect 4816 15200 4832 15264
rect 4896 15200 4912 15264
rect 4976 15200 4992 15264
rect 5056 15200 5064 15264
rect 4744 15046 5064 15200
rect 4744 14810 4786 15046
rect 5022 14810 5064 15046
rect 4744 14176 5064 14810
rect 4744 14112 4752 14176
rect 4816 14112 4832 14176
rect 4896 14112 4912 14176
rect 4976 14112 4992 14176
rect 5056 14112 5064 14176
rect 4744 13088 5064 14112
rect 4744 13024 4752 13088
rect 4816 13024 4832 13088
rect 4896 13024 4912 13088
rect 4976 13024 4992 13088
rect 5056 13024 5064 13088
rect 4744 12046 5064 13024
rect 4744 12000 4786 12046
rect 5022 12000 5064 12046
rect 4744 11936 4752 12000
rect 5056 11936 5064 12000
rect 4744 11810 4786 11936
rect 5022 11810 5064 11936
rect 4744 10912 5064 11810
rect 4744 10848 4752 10912
rect 4816 10848 4832 10912
rect 4896 10848 4912 10912
rect 4976 10848 4992 10912
rect 5056 10848 5064 10912
rect 4744 9824 5064 10848
rect 4744 9760 4752 9824
rect 4816 9760 4832 9824
rect 4896 9760 4912 9824
rect 4976 9760 4992 9824
rect 5056 9760 5064 9824
rect 4744 9046 5064 9760
rect 4744 8810 4786 9046
rect 5022 8810 5064 9046
rect 4744 8736 5064 8810
rect 4744 8672 4752 8736
rect 4816 8672 4832 8736
rect 4896 8672 4912 8736
rect 4976 8672 4992 8736
rect 5056 8672 5064 8736
rect 4744 7648 5064 8672
rect 4744 7584 4752 7648
rect 4816 7584 4832 7648
rect 4896 7584 4912 7648
rect 4976 7584 4992 7648
rect 5056 7584 5064 7648
rect 4744 6560 5064 7584
rect 4744 6496 4752 6560
rect 4816 6496 4832 6560
rect 4896 6496 4912 6560
rect 4976 6496 4992 6560
rect 5056 6496 5064 6560
rect 4744 6046 5064 6496
rect 4744 5810 4786 6046
rect 5022 5810 5064 6046
rect 4744 5472 5064 5810
rect 4744 5408 4752 5472
rect 4816 5408 4832 5472
rect 4896 5408 4912 5472
rect 4976 5408 4992 5472
rect 5056 5408 5064 5472
rect 4744 4384 5064 5408
rect 4744 4320 4752 4384
rect 4816 4320 4832 4384
rect 4896 4320 4912 4384
rect 4976 4320 4992 4384
rect 5056 4320 5064 4384
rect 4744 3296 5064 4320
rect 4744 3232 4752 3296
rect 4816 3232 4832 3296
rect 4896 3232 4912 3296
rect 4976 3232 4992 3296
rect 5056 3232 5064 3296
rect 4744 3046 5064 3232
rect 4744 2810 4786 3046
rect 5022 2810 5064 3046
rect 4744 2208 5064 2810
rect 4744 2144 4752 2208
rect 4816 2144 4832 2208
rect 4896 2144 4912 2208
rect 4976 2144 4992 2208
rect 5056 2144 5064 2208
rect 4744 2128 5064 2144
rect 6244 28864 6564 29424
rect 6244 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6412 28864
rect 6476 28800 6492 28864
rect 6556 28800 6564 28864
rect 6244 28546 6564 28800
rect 6244 28310 6286 28546
rect 6522 28310 6564 28546
rect 6244 27776 6564 28310
rect 6244 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6412 27776
rect 6476 27712 6492 27776
rect 6556 27712 6564 27776
rect 6244 26688 6564 27712
rect 6244 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6412 26688
rect 6476 26624 6492 26688
rect 6556 26624 6564 26688
rect 6244 25600 6564 26624
rect 6244 25536 6252 25600
rect 6316 25546 6332 25600
rect 6396 25546 6412 25600
rect 6476 25546 6492 25600
rect 6556 25536 6564 25600
rect 6244 25310 6286 25536
rect 6522 25310 6564 25536
rect 6244 24512 6564 25310
rect 6244 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6412 24512
rect 6476 24448 6492 24512
rect 6556 24448 6564 24512
rect 6244 23424 6564 24448
rect 6244 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6412 23424
rect 6476 23360 6492 23424
rect 6556 23360 6564 23424
rect 6244 22546 6564 23360
rect 6244 22336 6286 22546
rect 6522 22336 6564 22546
rect 6244 22272 6252 22336
rect 6316 22272 6332 22310
rect 6396 22272 6412 22310
rect 6476 22272 6492 22310
rect 6556 22272 6564 22336
rect 6244 21248 6564 22272
rect 6244 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6412 21248
rect 6476 21184 6492 21248
rect 6556 21184 6564 21248
rect 6244 20160 6564 21184
rect 6244 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6412 20160
rect 6476 20096 6492 20160
rect 6556 20096 6564 20160
rect 6244 19546 6564 20096
rect 6244 19310 6286 19546
rect 6522 19310 6564 19546
rect 6244 19072 6564 19310
rect 6244 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6412 19072
rect 6476 19008 6492 19072
rect 6556 19008 6564 19072
rect 6244 17984 6564 19008
rect 6244 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6412 17984
rect 6476 17920 6492 17984
rect 6556 17920 6564 17984
rect 6244 16896 6564 17920
rect 6244 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6412 16896
rect 6476 16832 6492 16896
rect 6556 16832 6564 16896
rect 6244 16546 6564 16832
rect 6244 16310 6286 16546
rect 6522 16310 6564 16546
rect 6244 15808 6564 16310
rect 6244 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6412 15808
rect 6476 15744 6492 15808
rect 6556 15744 6564 15808
rect 6244 14720 6564 15744
rect 6244 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6412 14720
rect 6476 14656 6492 14720
rect 6556 14656 6564 14720
rect 6244 13632 6564 14656
rect 6244 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6412 13632
rect 6476 13568 6492 13632
rect 6556 13568 6564 13632
rect 6244 13546 6564 13568
rect 6244 13310 6286 13546
rect 6522 13310 6564 13546
rect 6244 12544 6564 13310
rect 6244 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6412 12544
rect 6476 12480 6492 12544
rect 6556 12480 6564 12544
rect 6244 11456 6564 12480
rect 6244 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6412 11456
rect 6476 11392 6492 11456
rect 6556 11392 6564 11456
rect 6244 10546 6564 11392
rect 6244 10368 6286 10546
rect 6522 10368 6564 10546
rect 6244 10304 6252 10368
rect 6316 10304 6332 10310
rect 6396 10304 6412 10310
rect 6476 10304 6492 10310
rect 6556 10304 6564 10368
rect 6244 9280 6564 10304
rect 6244 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6412 9280
rect 6476 9216 6492 9280
rect 6556 9216 6564 9280
rect 6244 8192 6564 9216
rect 6244 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6412 8192
rect 6476 8128 6492 8192
rect 6556 8128 6564 8192
rect 6244 7546 6564 8128
rect 6244 7310 6286 7546
rect 6522 7310 6564 7546
rect 6244 7104 6564 7310
rect 6244 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6412 7104
rect 6476 7040 6492 7104
rect 6556 7040 6564 7104
rect 6244 6016 6564 7040
rect 6244 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6412 6016
rect 6476 5952 6492 6016
rect 6556 5952 6564 6016
rect 6244 4928 6564 5952
rect 6244 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6412 4928
rect 6476 4864 6492 4928
rect 6556 4864 6564 4928
rect 6244 4546 6564 4864
rect 6244 4310 6286 4546
rect 6522 4310 6564 4546
rect 6244 3840 6564 4310
rect 6244 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6412 3840
rect 6476 3776 6492 3840
rect 6556 3776 6564 3840
rect 6244 2752 6564 3776
rect 6244 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6412 2752
rect 6476 2688 6492 2752
rect 6556 2688 6564 2752
rect 6244 2128 6564 2688
rect 7744 29408 8064 29424
rect 7744 29344 7752 29408
rect 7816 29344 7832 29408
rect 7896 29344 7912 29408
rect 7976 29344 7992 29408
rect 8056 29344 8064 29408
rect 7744 28320 8064 29344
rect 7744 28256 7752 28320
rect 7816 28256 7832 28320
rect 7896 28256 7912 28320
rect 7976 28256 7992 28320
rect 8056 28256 8064 28320
rect 7744 27232 8064 28256
rect 7744 27168 7752 27232
rect 7816 27168 7832 27232
rect 7896 27168 7912 27232
rect 7976 27168 7992 27232
rect 8056 27168 8064 27232
rect 7744 27046 8064 27168
rect 7744 26810 7786 27046
rect 8022 26810 8064 27046
rect 7744 26144 8064 26810
rect 7744 26080 7752 26144
rect 7816 26080 7832 26144
rect 7896 26080 7912 26144
rect 7976 26080 7992 26144
rect 8056 26080 8064 26144
rect 7744 25056 8064 26080
rect 7744 24992 7752 25056
rect 7816 24992 7832 25056
rect 7896 24992 7912 25056
rect 7976 24992 7992 25056
rect 8056 24992 8064 25056
rect 7744 24046 8064 24992
rect 7744 23968 7786 24046
rect 8022 23968 8064 24046
rect 7744 23904 7752 23968
rect 8056 23904 8064 23968
rect 7744 23810 7786 23904
rect 8022 23810 8064 23904
rect 7744 22880 8064 23810
rect 7744 22816 7752 22880
rect 7816 22816 7832 22880
rect 7896 22816 7912 22880
rect 7976 22816 7992 22880
rect 8056 22816 8064 22880
rect 7744 21792 8064 22816
rect 7744 21728 7752 21792
rect 7816 21728 7832 21792
rect 7896 21728 7912 21792
rect 7976 21728 7992 21792
rect 8056 21728 8064 21792
rect 7744 21046 8064 21728
rect 7744 20810 7786 21046
rect 8022 20810 8064 21046
rect 7744 20704 8064 20810
rect 7744 20640 7752 20704
rect 7816 20640 7832 20704
rect 7896 20640 7912 20704
rect 7976 20640 7992 20704
rect 8056 20640 8064 20704
rect 7744 19616 8064 20640
rect 7744 19552 7752 19616
rect 7816 19552 7832 19616
rect 7896 19552 7912 19616
rect 7976 19552 7992 19616
rect 8056 19552 8064 19616
rect 7744 18528 8064 19552
rect 7744 18464 7752 18528
rect 7816 18464 7832 18528
rect 7896 18464 7912 18528
rect 7976 18464 7992 18528
rect 8056 18464 8064 18528
rect 7744 18046 8064 18464
rect 7744 17810 7786 18046
rect 8022 17810 8064 18046
rect 7744 17440 8064 17810
rect 7744 17376 7752 17440
rect 7816 17376 7832 17440
rect 7896 17376 7912 17440
rect 7976 17376 7992 17440
rect 8056 17376 8064 17440
rect 7744 16352 8064 17376
rect 7744 16288 7752 16352
rect 7816 16288 7832 16352
rect 7896 16288 7912 16352
rect 7976 16288 7992 16352
rect 8056 16288 8064 16352
rect 7744 15264 8064 16288
rect 7744 15200 7752 15264
rect 7816 15200 7832 15264
rect 7896 15200 7912 15264
rect 7976 15200 7992 15264
rect 8056 15200 8064 15264
rect 7744 15046 8064 15200
rect 7744 14810 7786 15046
rect 8022 14810 8064 15046
rect 7744 14176 8064 14810
rect 7744 14112 7752 14176
rect 7816 14112 7832 14176
rect 7896 14112 7912 14176
rect 7976 14112 7992 14176
rect 8056 14112 8064 14176
rect 7744 13088 8064 14112
rect 7744 13024 7752 13088
rect 7816 13024 7832 13088
rect 7896 13024 7912 13088
rect 7976 13024 7992 13088
rect 8056 13024 8064 13088
rect 7744 12046 8064 13024
rect 7744 12000 7786 12046
rect 8022 12000 8064 12046
rect 7744 11936 7752 12000
rect 8056 11936 8064 12000
rect 7744 11810 7786 11936
rect 8022 11810 8064 11936
rect 7744 10912 8064 11810
rect 7744 10848 7752 10912
rect 7816 10848 7832 10912
rect 7896 10848 7912 10912
rect 7976 10848 7992 10912
rect 8056 10848 8064 10912
rect 7744 9824 8064 10848
rect 7744 9760 7752 9824
rect 7816 9760 7832 9824
rect 7896 9760 7912 9824
rect 7976 9760 7992 9824
rect 8056 9760 8064 9824
rect 7744 9046 8064 9760
rect 7744 8810 7786 9046
rect 8022 8810 8064 9046
rect 7744 8736 8064 8810
rect 7744 8672 7752 8736
rect 7816 8672 7832 8736
rect 7896 8672 7912 8736
rect 7976 8672 7992 8736
rect 8056 8672 8064 8736
rect 7744 7648 8064 8672
rect 7744 7584 7752 7648
rect 7816 7584 7832 7648
rect 7896 7584 7912 7648
rect 7976 7584 7992 7648
rect 8056 7584 8064 7648
rect 7744 6560 8064 7584
rect 7744 6496 7752 6560
rect 7816 6496 7832 6560
rect 7896 6496 7912 6560
rect 7976 6496 7992 6560
rect 8056 6496 8064 6560
rect 7744 6046 8064 6496
rect 7744 5810 7786 6046
rect 8022 5810 8064 6046
rect 7744 5472 8064 5810
rect 7744 5408 7752 5472
rect 7816 5408 7832 5472
rect 7896 5408 7912 5472
rect 7976 5408 7992 5472
rect 8056 5408 8064 5472
rect 7744 4384 8064 5408
rect 7744 4320 7752 4384
rect 7816 4320 7832 4384
rect 7896 4320 7912 4384
rect 7976 4320 7992 4384
rect 8056 4320 8064 4384
rect 7744 3296 8064 4320
rect 7744 3232 7752 3296
rect 7816 3232 7832 3296
rect 7896 3232 7912 3296
rect 7976 3232 7992 3296
rect 8056 3232 8064 3296
rect 7744 3046 8064 3232
rect 7744 2810 7786 3046
rect 8022 2810 8064 3046
rect 7744 2208 8064 2810
rect 7744 2144 7752 2208
rect 7816 2144 7832 2208
rect 7896 2144 7912 2208
rect 7976 2144 7992 2208
rect 8056 2144 8064 2208
rect 7744 2128 8064 2144
rect 9244 28864 9564 29424
rect 9244 28800 9252 28864
rect 9316 28800 9332 28864
rect 9396 28800 9412 28864
rect 9476 28800 9492 28864
rect 9556 28800 9564 28864
rect 9244 28546 9564 28800
rect 9244 28310 9286 28546
rect 9522 28310 9564 28546
rect 9244 27776 9564 28310
rect 9244 27712 9252 27776
rect 9316 27712 9332 27776
rect 9396 27712 9412 27776
rect 9476 27712 9492 27776
rect 9556 27712 9564 27776
rect 9244 26688 9564 27712
rect 9244 26624 9252 26688
rect 9316 26624 9332 26688
rect 9396 26624 9412 26688
rect 9476 26624 9492 26688
rect 9556 26624 9564 26688
rect 9244 25600 9564 26624
rect 9244 25536 9252 25600
rect 9316 25546 9332 25600
rect 9396 25546 9412 25600
rect 9476 25546 9492 25600
rect 9556 25536 9564 25600
rect 9244 25310 9286 25536
rect 9522 25310 9564 25536
rect 9244 24512 9564 25310
rect 9244 24448 9252 24512
rect 9316 24448 9332 24512
rect 9396 24448 9412 24512
rect 9476 24448 9492 24512
rect 9556 24448 9564 24512
rect 9244 23424 9564 24448
rect 9244 23360 9252 23424
rect 9316 23360 9332 23424
rect 9396 23360 9412 23424
rect 9476 23360 9492 23424
rect 9556 23360 9564 23424
rect 9244 22546 9564 23360
rect 9244 22336 9286 22546
rect 9522 22336 9564 22546
rect 9244 22272 9252 22336
rect 9316 22272 9332 22310
rect 9396 22272 9412 22310
rect 9476 22272 9492 22310
rect 9556 22272 9564 22336
rect 9244 21248 9564 22272
rect 9244 21184 9252 21248
rect 9316 21184 9332 21248
rect 9396 21184 9412 21248
rect 9476 21184 9492 21248
rect 9556 21184 9564 21248
rect 9244 20160 9564 21184
rect 9244 20096 9252 20160
rect 9316 20096 9332 20160
rect 9396 20096 9412 20160
rect 9476 20096 9492 20160
rect 9556 20096 9564 20160
rect 9244 19546 9564 20096
rect 9244 19310 9286 19546
rect 9522 19310 9564 19546
rect 9244 19072 9564 19310
rect 9244 19008 9252 19072
rect 9316 19008 9332 19072
rect 9396 19008 9412 19072
rect 9476 19008 9492 19072
rect 9556 19008 9564 19072
rect 9244 17984 9564 19008
rect 9244 17920 9252 17984
rect 9316 17920 9332 17984
rect 9396 17920 9412 17984
rect 9476 17920 9492 17984
rect 9556 17920 9564 17984
rect 9244 16896 9564 17920
rect 9244 16832 9252 16896
rect 9316 16832 9332 16896
rect 9396 16832 9412 16896
rect 9476 16832 9492 16896
rect 9556 16832 9564 16896
rect 9244 16546 9564 16832
rect 9244 16310 9286 16546
rect 9522 16310 9564 16546
rect 9244 15808 9564 16310
rect 9244 15744 9252 15808
rect 9316 15744 9332 15808
rect 9396 15744 9412 15808
rect 9476 15744 9492 15808
rect 9556 15744 9564 15808
rect 9244 14720 9564 15744
rect 9244 14656 9252 14720
rect 9316 14656 9332 14720
rect 9396 14656 9412 14720
rect 9476 14656 9492 14720
rect 9556 14656 9564 14720
rect 9244 13632 9564 14656
rect 9244 13568 9252 13632
rect 9316 13568 9332 13632
rect 9396 13568 9412 13632
rect 9476 13568 9492 13632
rect 9556 13568 9564 13632
rect 9244 13546 9564 13568
rect 9244 13310 9286 13546
rect 9522 13310 9564 13546
rect 9244 12544 9564 13310
rect 9244 12480 9252 12544
rect 9316 12480 9332 12544
rect 9396 12480 9412 12544
rect 9476 12480 9492 12544
rect 9556 12480 9564 12544
rect 9244 11456 9564 12480
rect 9244 11392 9252 11456
rect 9316 11392 9332 11456
rect 9396 11392 9412 11456
rect 9476 11392 9492 11456
rect 9556 11392 9564 11456
rect 9244 10546 9564 11392
rect 9244 10368 9286 10546
rect 9522 10368 9564 10546
rect 9244 10304 9252 10368
rect 9316 10304 9332 10310
rect 9396 10304 9412 10310
rect 9476 10304 9492 10310
rect 9556 10304 9564 10368
rect 9244 9280 9564 10304
rect 9244 9216 9252 9280
rect 9316 9216 9332 9280
rect 9396 9216 9412 9280
rect 9476 9216 9492 9280
rect 9556 9216 9564 9280
rect 9244 8192 9564 9216
rect 9244 8128 9252 8192
rect 9316 8128 9332 8192
rect 9396 8128 9412 8192
rect 9476 8128 9492 8192
rect 9556 8128 9564 8192
rect 9244 7546 9564 8128
rect 9244 7310 9286 7546
rect 9522 7310 9564 7546
rect 9244 7104 9564 7310
rect 9244 7040 9252 7104
rect 9316 7040 9332 7104
rect 9396 7040 9412 7104
rect 9476 7040 9492 7104
rect 9556 7040 9564 7104
rect 9244 6016 9564 7040
rect 9244 5952 9252 6016
rect 9316 5952 9332 6016
rect 9396 5952 9412 6016
rect 9476 5952 9492 6016
rect 9556 5952 9564 6016
rect 9244 4928 9564 5952
rect 9244 4864 9252 4928
rect 9316 4864 9332 4928
rect 9396 4864 9412 4928
rect 9476 4864 9492 4928
rect 9556 4864 9564 4928
rect 9244 4546 9564 4864
rect 9244 4310 9286 4546
rect 9522 4310 9564 4546
rect 9244 3840 9564 4310
rect 9244 3776 9252 3840
rect 9316 3776 9332 3840
rect 9396 3776 9412 3840
rect 9476 3776 9492 3840
rect 9556 3776 9564 3840
rect 9244 2752 9564 3776
rect 9244 2688 9252 2752
rect 9316 2688 9332 2752
rect 9396 2688 9412 2752
rect 9476 2688 9492 2752
rect 9556 2688 9564 2752
rect 9244 2128 9564 2688
rect 10744 29408 11064 29424
rect 10744 29344 10752 29408
rect 10816 29344 10832 29408
rect 10896 29344 10912 29408
rect 10976 29344 10992 29408
rect 11056 29344 11064 29408
rect 10744 28320 11064 29344
rect 10744 28256 10752 28320
rect 10816 28256 10832 28320
rect 10896 28256 10912 28320
rect 10976 28256 10992 28320
rect 11056 28256 11064 28320
rect 10744 27232 11064 28256
rect 10744 27168 10752 27232
rect 10816 27168 10832 27232
rect 10896 27168 10912 27232
rect 10976 27168 10992 27232
rect 11056 27168 11064 27232
rect 10744 27046 11064 27168
rect 10744 26810 10786 27046
rect 11022 26810 11064 27046
rect 10744 26144 11064 26810
rect 10744 26080 10752 26144
rect 10816 26080 10832 26144
rect 10896 26080 10912 26144
rect 10976 26080 10992 26144
rect 11056 26080 11064 26144
rect 10744 25056 11064 26080
rect 10744 24992 10752 25056
rect 10816 24992 10832 25056
rect 10896 24992 10912 25056
rect 10976 24992 10992 25056
rect 11056 24992 11064 25056
rect 10744 24046 11064 24992
rect 10744 23968 10786 24046
rect 11022 23968 11064 24046
rect 10744 23904 10752 23968
rect 11056 23904 11064 23968
rect 10744 23810 10786 23904
rect 11022 23810 11064 23904
rect 10744 22880 11064 23810
rect 10744 22816 10752 22880
rect 10816 22816 10832 22880
rect 10896 22816 10912 22880
rect 10976 22816 10992 22880
rect 11056 22816 11064 22880
rect 10744 21792 11064 22816
rect 10744 21728 10752 21792
rect 10816 21728 10832 21792
rect 10896 21728 10912 21792
rect 10976 21728 10992 21792
rect 11056 21728 11064 21792
rect 10744 21046 11064 21728
rect 10744 20810 10786 21046
rect 11022 20810 11064 21046
rect 10744 20704 11064 20810
rect 10744 20640 10752 20704
rect 10816 20640 10832 20704
rect 10896 20640 10912 20704
rect 10976 20640 10992 20704
rect 11056 20640 11064 20704
rect 10744 19616 11064 20640
rect 10744 19552 10752 19616
rect 10816 19552 10832 19616
rect 10896 19552 10912 19616
rect 10976 19552 10992 19616
rect 11056 19552 11064 19616
rect 10744 18528 11064 19552
rect 10744 18464 10752 18528
rect 10816 18464 10832 18528
rect 10896 18464 10912 18528
rect 10976 18464 10992 18528
rect 11056 18464 11064 18528
rect 10744 18046 11064 18464
rect 10744 17810 10786 18046
rect 11022 17810 11064 18046
rect 10744 17440 11064 17810
rect 10744 17376 10752 17440
rect 10816 17376 10832 17440
rect 10896 17376 10912 17440
rect 10976 17376 10992 17440
rect 11056 17376 11064 17440
rect 10744 16352 11064 17376
rect 10744 16288 10752 16352
rect 10816 16288 10832 16352
rect 10896 16288 10912 16352
rect 10976 16288 10992 16352
rect 11056 16288 11064 16352
rect 10744 15264 11064 16288
rect 10744 15200 10752 15264
rect 10816 15200 10832 15264
rect 10896 15200 10912 15264
rect 10976 15200 10992 15264
rect 11056 15200 11064 15264
rect 10744 15046 11064 15200
rect 10744 14810 10786 15046
rect 11022 14810 11064 15046
rect 10744 14176 11064 14810
rect 10744 14112 10752 14176
rect 10816 14112 10832 14176
rect 10896 14112 10912 14176
rect 10976 14112 10992 14176
rect 11056 14112 11064 14176
rect 10744 13088 11064 14112
rect 10744 13024 10752 13088
rect 10816 13024 10832 13088
rect 10896 13024 10912 13088
rect 10976 13024 10992 13088
rect 11056 13024 11064 13088
rect 10744 12046 11064 13024
rect 10744 12000 10786 12046
rect 11022 12000 11064 12046
rect 10744 11936 10752 12000
rect 11056 11936 11064 12000
rect 10744 11810 10786 11936
rect 11022 11810 11064 11936
rect 10744 10912 11064 11810
rect 10744 10848 10752 10912
rect 10816 10848 10832 10912
rect 10896 10848 10912 10912
rect 10976 10848 10992 10912
rect 11056 10848 11064 10912
rect 10744 9824 11064 10848
rect 10744 9760 10752 9824
rect 10816 9760 10832 9824
rect 10896 9760 10912 9824
rect 10976 9760 10992 9824
rect 11056 9760 11064 9824
rect 10744 9046 11064 9760
rect 10744 8810 10786 9046
rect 11022 8810 11064 9046
rect 10744 8736 11064 8810
rect 10744 8672 10752 8736
rect 10816 8672 10832 8736
rect 10896 8672 10912 8736
rect 10976 8672 10992 8736
rect 11056 8672 11064 8736
rect 10744 7648 11064 8672
rect 10744 7584 10752 7648
rect 10816 7584 10832 7648
rect 10896 7584 10912 7648
rect 10976 7584 10992 7648
rect 11056 7584 11064 7648
rect 10744 6560 11064 7584
rect 10744 6496 10752 6560
rect 10816 6496 10832 6560
rect 10896 6496 10912 6560
rect 10976 6496 10992 6560
rect 11056 6496 11064 6560
rect 10744 6046 11064 6496
rect 10744 5810 10786 6046
rect 11022 5810 11064 6046
rect 10744 5472 11064 5810
rect 10744 5408 10752 5472
rect 10816 5408 10832 5472
rect 10896 5408 10912 5472
rect 10976 5408 10992 5472
rect 11056 5408 11064 5472
rect 10744 4384 11064 5408
rect 10744 4320 10752 4384
rect 10816 4320 10832 4384
rect 10896 4320 10912 4384
rect 10976 4320 10992 4384
rect 11056 4320 11064 4384
rect 10744 3296 11064 4320
rect 10744 3232 10752 3296
rect 10816 3232 10832 3296
rect 10896 3232 10912 3296
rect 10976 3232 10992 3296
rect 11056 3232 11064 3296
rect 10744 3046 11064 3232
rect 10744 2810 10786 3046
rect 11022 2810 11064 3046
rect 10744 2208 11064 2810
rect 10744 2144 10752 2208
rect 10816 2144 10832 2208
rect 10896 2144 10912 2208
rect 10976 2144 10992 2208
rect 11056 2144 11064 2208
rect 10744 2128 11064 2144
rect 12244 28864 12564 29424
rect 12244 28800 12252 28864
rect 12316 28800 12332 28864
rect 12396 28800 12412 28864
rect 12476 28800 12492 28864
rect 12556 28800 12564 28864
rect 12244 28546 12564 28800
rect 12244 28310 12286 28546
rect 12522 28310 12564 28546
rect 12244 27776 12564 28310
rect 12244 27712 12252 27776
rect 12316 27712 12332 27776
rect 12396 27712 12412 27776
rect 12476 27712 12492 27776
rect 12556 27712 12564 27776
rect 12244 26688 12564 27712
rect 12244 26624 12252 26688
rect 12316 26624 12332 26688
rect 12396 26624 12412 26688
rect 12476 26624 12492 26688
rect 12556 26624 12564 26688
rect 12244 25600 12564 26624
rect 12244 25536 12252 25600
rect 12316 25546 12332 25600
rect 12396 25546 12412 25600
rect 12476 25546 12492 25600
rect 12556 25536 12564 25600
rect 12244 25310 12286 25536
rect 12522 25310 12564 25536
rect 12244 24512 12564 25310
rect 12244 24448 12252 24512
rect 12316 24448 12332 24512
rect 12396 24448 12412 24512
rect 12476 24448 12492 24512
rect 12556 24448 12564 24512
rect 12244 23424 12564 24448
rect 12244 23360 12252 23424
rect 12316 23360 12332 23424
rect 12396 23360 12412 23424
rect 12476 23360 12492 23424
rect 12556 23360 12564 23424
rect 12244 22546 12564 23360
rect 12244 22336 12286 22546
rect 12522 22336 12564 22546
rect 12244 22272 12252 22336
rect 12316 22272 12332 22310
rect 12396 22272 12412 22310
rect 12476 22272 12492 22310
rect 12556 22272 12564 22336
rect 12244 21248 12564 22272
rect 12244 21184 12252 21248
rect 12316 21184 12332 21248
rect 12396 21184 12412 21248
rect 12476 21184 12492 21248
rect 12556 21184 12564 21248
rect 12244 20160 12564 21184
rect 12244 20096 12252 20160
rect 12316 20096 12332 20160
rect 12396 20096 12412 20160
rect 12476 20096 12492 20160
rect 12556 20096 12564 20160
rect 12244 19546 12564 20096
rect 12244 19310 12286 19546
rect 12522 19310 12564 19546
rect 12244 19072 12564 19310
rect 12244 19008 12252 19072
rect 12316 19008 12332 19072
rect 12396 19008 12412 19072
rect 12476 19008 12492 19072
rect 12556 19008 12564 19072
rect 12244 17984 12564 19008
rect 12244 17920 12252 17984
rect 12316 17920 12332 17984
rect 12396 17920 12412 17984
rect 12476 17920 12492 17984
rect 12556 17920 12564 17984
rect 12244 16896 12564 17920
rect 12244 16832 12252 16896
rect 12316 16832 12332 16896
rect 12396 16832 12412 16896
rect 12476 16832 12492 16896
rect 12556 16832 12564 16896
rect 12244 16546 12564 16832
rect 12244 16310 12286 16546
rect 12522 16310 12564 16546
rect 12244 15808 12564 16310
rect 12244 15744 12252 15808
rect 12316 15744 12332 15808
rect 12396 15744 12412 15808
rect 12476 15744 12492 15808
rect 12556 15744 12564 15808
rect 12244 14720 12564 15744
rect 12244 14656 12252 14720
rect 12316 14656 12332 14720
rect 12396 14656 12412 14720
rect 12476 14656 12492 14720
rect 12556 14656 12564 14720
rect 12244 13632 12564 14656
rect 12244 13568 12252 13632
rect 12316 13568 12332 13632
rect 12396 13568 12412 13632
rect 12476 13568 12492 13632
rect 12556 13568 12564 13632
rect 12244 13546 12564 13568
rect 12244 13310 12286 13546
rect 12522 13310 12564 13546
rect 12244 12544 12564 13310
rect 12244 12480 12252 12544
rect 12316 12480 12332 12544
rect 12396 12480 12412 12544
rect 12476 12480 12492 12544
rect 12556 12480 12564 12544
rect 12244 11456 12564 12480
rect 12244 11392 12252 11456
rect 12316 11392 12332 11456
rect 12396 11392 12412 11456
rect 12476 11392 12492 11456
rect 12556 11392 12564 11456
rect 12244 10546 12564 11392
rect 12244 10368 12286 10546
rect 12522 10368 12564 10546
rect 12244 10304 12252 10368
rect 12316 10304 12332 10310
rect 12396 10304 12412 10310
rect 12476 10304 12492 10310
rect 12556 10304 12564 10368
rect 12244 9280 12564 10304
rect 12244 9216 12252 9280
rect 12316 9216 12332 9280
rect 12396 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12564 9280
rect 12244 8192 12564 9216
rect 12244 8128 12252 8192
rect 12316 8128 12332 8192
rect 12396 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12564 8192
rect 12244 7546 12564 8128
rect 12244 7310 12286 7546
rect 12522 7310 12564 7546
rect 12244 7104 12564 7310
rect 12244 7040 12252 7104
rect 12316 7040 12332 7104
rect 12396 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12564 7104
rect 12244 6016 12564 7040
rect 12244 5952 12252 6016
rect 12316 5952 12332 6016
rect 12396 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12564 6016
rect 12244 4928 12564 5952
rect 12244 4864 12252 4928
rect 12316 4864 12332 4928
rect 12396 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12564 4928
rect 12244 4546 12564 4864
rect 12244 4310 12286 4546
rect 12522 4310 12564 4546
rect 12244 3840 12564 4310
rect 12244 3776 12252 3840
rect 12316 3776 12332 3840
rect 12396 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12564 3840
rect 12244 2752 12564 3776
rect 12244 2688 12252 2752
rect 12316 2688 12332 2752
rect 12396 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12564 2752
rect 12244 2128 12564 2688
rect 13744 29408 14064 29424
rect 13744 29344 13752 29408
rect 13816 29344 13832 29408
rect 13896 29344 13912 29408
rect 13976 29344 13992 29408
rect 14056 29344 14064 29408
rect 13744 28320 14064 29344
rect 13744 28256 13752 28320
rect 13816 28256 13832 28320
rect 13896 28256 13912 28320
rect 13976 28256 13992 28320
rect 14056 28256 14064 28320
rect 13744 27232 14064 28256
rect 13744 27168 13752 27232
rect 13816 27168 13832 27232
rect 13896 27168 13912 27232
rect 13976 27168 13992 27232
rect 14056 27168 14064 27232
rect 13744 27046 14064 27168
rect 13744 26810 13786 27046
rect 14022 26810 14064 27046
rect 13744 26144 14064 26810
rect 13744 26080 13752 26144
rect 13816 26080 13832 26144
rect 13896 26080 13912 26144
rect 13976 26080 13992 26144
rect 14056 26080 14064 26144
rect 13744 25056 14064 26080
rect 13744 24992 13752 25056
rect 13816 24992 13832 25056
rect 13896 24992 13912 25056
rect 13976 24992 13992 25056
rect 14056 24992 14064 25056
rect 13744 24046 14064 24992
rect 13744 23968 13786 24046
rect 14022 23968 14064 24046
rect 13744 23904 13752 23968
rect 14056 23904 14064 23968
rect 13744 23810 13786 23904
rect 14022 23810 14064 23904
rect 13744 22880 14064 23810
rect 13744 22816 13752 22880
rect 13816 22816 13832 22880
rect 13896 22816 13912 22880
rect 13976 22816 13992 22880
rect 14056 22816 14064 22880
rect 13744 21792 14064 22816
rect 13744 21728 13752 21792
rect 13816 21728 13832 21792
rect 13896 21728 13912 21792
rect 13976 21728 13992 21792
rect 14056 21728 14064 21792
rect 13744 21046 14064 21728
rect 13744 20810 13786 21046
rect 14022 20810 14064 21046
rect 13744 20704 14064 20810
rect 13744 20640 13752 20704
rect 13816 20640 13832 20704
rect 13896 20640 13912 20704
rect 13976 20640 13992 20704
rect 14056 20640 14064 20704
rect 13744 19616 14064 20640
rect 13744 19552 13752 19616
rect 13816 19552 13832 19616
rect 13896 19552 13912 19616
rect 13976 19552 13992 19616
rect 14056 19552 14064 19616
rect 13744 18528 14064 19552
rect 13744 18464 13752 18528
rect 13816 18464 13832 18528
rect 13896 18464 13912 18528
rect 13976 18464 13992 18528
rect 14056 18464 14064 18528
rect 13744 18046 14064 18464
rect 13744 17810 13786 18046
rect 14022 17810 14064 18046
rect 13744 17440 14064 17810
rect 13744 17376 13752 17440
rect 13816 17376 13832 17440
rect 13896 17376 13912 17440
rect 13976 17376 13992 17440
rect 14056 17376 14064 17440
rect 13744 16352 14064 17376
rect 13744 16288 13752 16352
rect 13816 16288 13832 16352
rect 13896 16288 13912 16352
rect 13976 16288 13992 16352
rect 14056 16288 14064 16352
rect 13744 15264 14064 16288
rect 13744 15200 13752 15264
rect 13816 15200 13832 15264
rect 13896 15200 13912 15264
rect 13976 15200 13992 15264
rect 14056 15200 14064 15264
rect 13744 15046 14064 15200
rect 13744 14810 13786 15046
rect 14022 14810 14064 15046
rect 13744 14176 14064 14810
rect 13744 14112 13752 14176
rect 13816 14112 13832 14176
rect 13896 14112 13912 14176
rect 13976 14112 13992 14176
rect 14056 14112 14064 14176
rect 13744 13088 14064 14112
rect 13744 13024 13752 13088
rect 13816 13024 13832 13088
rect 13896 13024 13912 13088
rect 13976 13024 13992 13088
rect 14056 13024 14064 13088
rect 13744 12046 14064 13024
rect 13744 12000 13786 12046
rect 14022 12000 14064 12046
rect 13744 11936 13752 12000
rect 14056 11936 14064 12000
rect 13744 11810 13786 11936
rect 14022 11810 14064 11936
rect 13744 10912 14064 11810
rect 13744 10848 13752 10912
rect 13816 10848 13832 10912
rect 13896 10848 13912 10912
rect 13976 10848 13992 10912
rect 14056 10848 14064 10912
rect 13744 9824 14064 10848
rect 13744 9760 13752 9824
rect 13816 9760 13832 9824
rect 13896 9760 13912 9824
rect 13976 9760 13992 9824
rect 14056 9760 14064 9824
rect 13744 9046 14064 9760
rect 13744 8810 13786 9046
rect 14022 8810 14064 9046
rect 13744 8736 14064 8810
rect 13744 8672 13752 8736
rect 13816 8672 13832 8736
rect 13896 8672 13912 8736
rect 13976 8672 13992 8736
rect 14056 8672 14064 8736
rect 13744 7648 14064 8672
rect 13744 7584 13752 7648
rect 13816 7584 13832 7648
rect 13896 7584 13912 7648
rect 13976 7584 13992 7648
rect 14056 7584 14064 7648
rect 13744 6560 14064 7584
rect 13744 6496 13752 6560
rect 13816 6496 13832 6560
rect 13896 6496 13912 6560
rect 13976 6496 13992 6560
rect 14056 6496 14064 6560
rect 13744 6046 14064 6496
rect 13744 5810 13786 6046
rect 14022 5810 14064 6046
rect 13744 5472 14064 5810
rect 13744 5408 13752 5472
rect 13816 5408 13832 5472
rect 13896 5408 13912 5472
rect 13976 5408 13992 5472
rect 14056 5408 14064 5472
rect 13744 4384 14064 5408
rect 13744 4320 13752 4384
rect 13816 4320 13832 4384
rect 13896 4320 13912 4384
rect 13976 4320 13992 4384
rect 14056 4320 14064 4384
rect 13744 3296 14064 4320
rect 13744 3232 13752 3296
rect 13816 3232 13832 3296
rect 13896 3232 13912 3296
rect 13976 3232 13992 3296
rect 14056 3232 14064 3296
rect 13744 3046 14064 3232
rect 13744 2810 13786 3046
rect 14022 2810 14064 3046
rect 13744 2208 14064 2810
rect 13744 2144 13752 2208
rect 13816 2144 13832 2208
rect 13896 2144 13912 2208
rect 13976 2144 13992 2208
rect 14056 2144 14064 2208
rect 13744 2128 14064 2144
rect 15244 28864 15564 29424
rect 15244 28800 15252 28864
rect 15316 28800 15332 28864
rect 15396 28800 15412 28864
rect 15476 28800 15492 28864
rect 15556 28800 15564 28864
rect 15244 28546 15564 28800
rect 15244 28310 15286 28546
rect 15522 28310 15564 28546
rect 15244 27776 15564 28310
rect 15244 27712 15252 27776
rect 15316 27712 15332 27776
rect 15396 27712 15412 27776
rect 15476 27712 15492 27776
rect 15556 27712 15564 27776
rect 15244 26688 15564 27712
rect 15244 26624 15252 26688
rect 15316 26624 15332 26688
rect 15396 26624 15412 26688
rect 15476 26624 15492 26688
rect 15556 26624 15564 26688
rect 15244 25600 15564 26624
rect 15244 25536 15252 25600
rect 15316 25546 15332 25600
rect 15396 25546 15412 25600
rect 15476 25546 15492 25600
rect 15556 25536 15564 25600
rect 15244 25310 15286 25536
rect 15522 25310 15564 25536
rect 15244 24512 15564 25310
rect 15244 24448 15252 24512
rect 15316 24448 15332 24512
rect 15396 24448 15412 24512
rect 15476 24448 15492 24512
rect 15556 24448 15564 24512
rect 15244 23424 15564 24448
rect 15244 23360 15252 23424
rect 15316 23360 15332 23424
rect 15396 23360 15412 23424
rect 15476 23360 15492 23424
rect 15556 23360 15564 23424
rect 15244 22546 15564 23360
rect 15244 22336 15286 22546
rect 15522 22336 15564 22546
rect 15244 22272 15252 22336
rect 15316 22272 15332 22310
rect 15396 22272 15412 22310
rect 15476 22272 15492 22310
rect 15556 22272 15564 22336
rect 15244 21248 15564 22272
rect 15244 21184 15252 21248
rect 15316 21184 15332 21248
rect 15396 21184 15412 21248
rect 15476 21184 15492 21248
rect 15556 21184 15564 21248
rect 15244 20160 15564 21184
rect 15244 20096 15252 20160
rect 15316 20096 15332 20160
rect 15396 20096 15412 20160
rect 15476 20096 15492 20160
rect 15556 20096 15564 20160
rect 15244 19546 15564 20096
rect 15244 19310 15286 19546
rect 15522 19310 15564 19546
rect 15244 19072 15564 19310
rect 15244 19008 15252 19072
rect 15316 19008 15332 19072
rect 15396 19008 15412 19072
rect 15476 19008 15492 19072
rect 15556 19008 15564 19072
rect 15244 17984 15564 19008
rect 15244 17920 15252 17984
rect 15316 17920 15332 17984
rect 15396 17920 15412 17984
rect 15476 17920 15492 17984
rect 15556 17920 15564 17984
rect 15244 16896 15564 17920
rect 15244 16832 15252 16896
rect 15316 16832 15332 16896
rect 15396 16832 15412 16896
rect 15476 16832 15492 16896
rect 15556 16832 15564 16896
rect 15244 16546 15564 16832
rect 15244 16310 15286 16546
rect 15522 16310 15564 16546
rect 15244 15808 15564 16310
rect 15244 15744 15252 15808
rect 15316 15744 15332 15808
rect 15396 15744 15412 15808
rect 15476 15744 15492 15808
rect 15556 15744 15564 15808
rect 15244 14720 15564 15744
rect 15244 14656 15252 14720
rect 15316 14656 15332 14720
rect 15396 14656 15412 14720
rect 15476 14656 15492 14720
rect 15556 14656 15564 14720
rect 15244 13632 15564 14656
rect 15244 13568 15252 13632
rect 15316 13568 15332 13632
rect 15396 13568 15412 13632
rect 15476 13568 15492 13632
rect 15556 13568 15564 13632
rect 15244 13546 15564 13568
rect 15244 13310 15286 13546
rect 15522 13310 15564 13546
rect 15244 12544 15564 13310
rect 15244 12480 15252 12544
rect 15316 12480 15332 12544
rect 15396 12480 15412 12544
rect 15476 12480 15492 12544
rect 15556 12480 15564 12544
rect 15244 11456 15564 12480
rect 15244 11392 15252 11456
rect 15316 11392 15332 11456
rect 15396 11392 15412 11456
rect 15476 11392 15492 11456
rect 15556 11392 15564 11456
rect 15244 10546 15564 11392
rect 15244 10368 15286 10546
rect 15522 10368 15564 10546
rect 15244 10304 15252 10368
rect 15316 10304 15332 10310
rect 15396 10304 15412 10310
rect 15476 10304 15492 10310
rect 15556 10304 15564 10368
rect 15244 9280 15564 10304
rect 15244 9216 15252 9280
rect 15316 9216 15332 9280
rect 15396 9216 15412 9280
rect 15476 9216 15492 9280
rect 15556 9216 15564 9280
rect 15244 8192 15564 9216
rect 15244 8128 15252 8192
rect 15316 8128 15332 8192
rect 15396 8128 15412 8192
rect 15476 8128 15492 8192
rect 15556 8128 15564 8192
rect 15244 7546 15564 8128
rect 15244 7310 15286 7546
rect 15522 7310 15564 7546
rect 15244 7104 15564 7310
rect 15244 7040 15252 7104
rect 15316 7040 15332 7104
rect 15396 7040 15412 7104
rect 15476 7040 15492 7104
rect 15556 7040 15564 7104
rect 15244 6016 15564 7040
rect 15244 5952 15252 6016
rect 15316 5952 15332 6016
rect 15396 5952 15412 6016
rect 15476 5952 15492 6016
rect 15556 5952 15564 6016
rect 15244 4928 15564 5952
rect 15244 4864 15252 4928
rect 15316 4864 15332 4928
rect 15396 4864 15412 4928
rect 15476 4864 15492 4928
rect 15556 4864 15564 4928
rect 15244 4546 15564 4864
rect 15244 4310 15286 4546
rect 15522 4310 15564 4546
rect 15244 3840 15564 4310
rect 15244 3776 15252 3840
rect 15316 3776 15332 3840
rect 15396 3776 15412 3840
rect 15476 3776 15492 3840
rect 15556 3776 15564 3840
rect 15244 2752 15564 3776
rect 15244 2688 15252 2752
rect 15316 2688 15332 2752
rect 15396 2688 15412 2752
rect 15476 2688 15492 2752
rect 15556 2688 15564 2752
rect 15244 2128 15564 2688
rect 16744 29408 17064 29424
rect 16744 29344 16752 29408
rect 16816 29344 16832 29408
rect 16896 29344 16912 29408
rect 16976 29344 16992 29408
rect 17056 29344 17064 29408
rect 16744 28320 17064 29344
rect 16744 28256 16752 28320
rect 16816 28256 16832 28320
rect 16896 28256 16912 28320
rect 16976 28256 16992 28320
rect 17056 28256 17064 28320
rect 16744 27232 17064 28256
rect 16744 27168 16752 27232
rect 16816 27168 16832 27232
rect 16896 27168 16912 27232
rect 16976 27168 16992 27232
rect 17056 27168 17064 27232
rect 16744 27046 17064 27168
rect 16744 26810 16786 27046
rect 17022 26810 17064 27046
rect 16744 26144 17064 26810
rect 16744 26080 16752 26144
rect 16816 26080 16832 26144
rect 16896 26080 16912 26144
rect 16976 26080 16992 26144
rect 17056 26080 17064 26144
rect 16744 25056 17064 26080
rect 16744 24992 16752 25056
rect 16816 24992 16832 25056
rect 16896 24992 16912 25056
rect 16976 24992 16992 25056
rect 17056 24992 17064 25056
rect 16744 24046 17064 24992
rect 16744 23968 16786 24046
rect 17022 23968 17064 24046
rect 16744 23904 16752 23968
rect 17056 23904 17064 23968
rect 16744 23810 16786 23904
rect 17022 23810 17064 23904
rect 16744 22880 17064 23810
rect 16744 22816 16752 22880
rect 16816 22816 16832 22880
rect 16896 22816 16912 22880
rect 16976 22816 16992 22880
rect 17056 22816 17064 22880
rect 16744 21792 17064 22816
rect 16744 21728 16752 21792
rect 16816 21728 16832 21792
rect 16896 21728 16912 21792
rect 16976 21728 16992 21792
rect 17056 21728 17064 21792
rect 16744 21046 17064 21728
rect 16744 20810 16786 21046
rect 17022 20810 17064 21046
rect 16744 20704 17064 20810
rect 16744 20640 16752 20704
rect 16816 20640 16832 20704
rect 16896 20640 16912 20704
rect 16976 20640 16992 20704
rect 17056 20640 17064 20704
rect 16744 19616 17064 20640
rect 16744 19552 16752 19616
rect 16816 19552 16832 19616
rect 16896 19552 16912 19616
rect 16976 19552 16992 19616
rect 17056 19552 17064 19616
rect 16744 18528 17064 19552
rect 16744 18464 16752 18528
rect 16816 18464 16832 18528
rect 16896 18464 16912 18528
rect 16976 18464 16992 18528
rect 17056 18464 17064 18528
rect 16744 18046 17064 18464
rect 16744 17810 16786 18046
rect 17022 17810 17064 18046
rect 16744 17440 17064 17810
rect 16744 17376 16752 17440
rect 16816 17376 16832 17440
rect 16896 17376 16912 17440
rect 16976 17376 16992 17440
rect 17056 17376 17064 17440
rect 16744 16352 17064 17376
rect 16744 16288 16752 16352
rect 16816 16288 16832 16352
rect 16896 16288 16912 16352
rect 16976 16288 16992 16352
rect 17056 16288 17064 16352
rect 16744 15264 17064 16288
rect 16744 15200 16752 15264
rect 16816 15200 16832 15264
rect 16896 15200 16912 15264
rect 16976 15200 16992 15264
rect 17056 15200 17064 15264
rect 16744 15046 17064 15200
rect 16744 14810 16786 15046
rect 17022 14810 17064 15046
rect 16744 14176 17064 14810
rect 16744 14112 16752 14176
rect 16816 14112 16832 14176
rect 16896 14112 16912 14176
rect 16976 14112 16992 14176
rect 17056 14112 17064 14176
rect 16744 13088 17064 14112
rect 16744 13024 16752 13088
rect 16816 13024 16832 13088
rect 16896 13024 16912 13088
rect 16976 13024 16992 13088
rect 17056 13024 17064 13088
rect 16744 12046 17064 13024
rect 16744 12000 16786 12046
rect 17022 12000 17064 12046
rect 16744 11936 16752 12000
rect 17056 11936 17064 12000
rect 16744 11810 16786 11936
rect 17022 11810 17064 11936
rect 16744 10912 17064 11810
rect 16744 10848 16752 10912
rect 16816 10848 16832 10912
rect 16896 10848 16912 10912
rect 16976 10848 16992 10912
rect 17056 10848 17064 10912
rect 16744 9824 17064 10848
rect 16744 9760 16752 9824
rect 16816 9760 16832 9824
rect 16896 9760 16912 9824
rect 16976 9760 16992 9824
rect 17056 9760 17064 9824
rect 16744 9046 17064 9760
rect 16744 8810 16786 9046
rect 17022 8810 17064 9046
rect 16744 8736 17064 8810
rect 16744 8672 16752 8736
rect 16816 8672 16832 8736
rect 16896 8672 16912 8736
rect 16976 8672 16992 8736
rect 17056 8672 17064 8736
rect 16744 7648 17064 8672
rect 16744 7584 16752 7648
rect 16816 7584 16832 7648
rect 16896 7584 16912 7648
rect 16976 7584 16992 7648
rect 17056 7584 17064 7648
rect 16744 6560 17064 7584
rect 16744 6496 16752 6560
rect 16816 6496 16832 6560
rect 16896 6496 16912 6560
rect 16976 6496 16992 6560
rect 17056 6496 17064 6560
rect 16744 6046 17064 6496
rect 16744 5810 16786 6046
rect 17022 5810 17064 6046
rect 16744 5472 17064 5810
rect 16744 5408 16752 5472
rect 16816 5408 16832 5472
rect 16896 5408 16912 5472
rect 16976 5408 16992 5472
rect 17056 5408 17064 5472
rect 16744 4384 17064 5408
rect 16744 4320 16752 4384
rect 16816 4320 16832 4384
rect 16896 4320 16912 4384
rect 16976 4320 16992 4384
rect 17056 4320 17064 4384
rect 16744 3296 17064 4320
rect 16744 3232 16752 3296
rect 16816 3232 16832 3296
rect 16896 3232 16912 3296
rect 16976 3232 16992 3296
rect 17056 3232 17064 3296
rect 16744 3046 17064 3232
rect 16744 2810 16786 3046
rect 17022 2810 17064 3046
rect 16744 2208 17064 2810
rect 16744 2144 16752 2208
rect 16816 2144 16832 2208
rect 16896 2144 16912 2208
rect 16976 2144 16992 2208
rect 17056 2144 17064 2208
rect 16744 2128 17064 2144
rect 18244 28864 18564 29424
rect 18244 28800 18252 28864
rect 18316 28800 18332 28864
rect 18396 28800 18412 28864
rect 18476 28800 18492 28864
rect 18556 28800 18564 28864
rect 18244 28546 18564 28800
rect 18244 28310 18286 28546
rect 18522 28310 18564 28546
rect 18244 27776 18564 28310
rect 18244 27712 18252 27776
rect 18316 27712 18332 27776
rect 18396 27712 18412 27776
rect 18476 27712 18492 27776
rect 18556 27712 18564 27776
rect 18244 26688 18564 27712
rect 18244 26624 18252 26688
rect 18316 26624 18332 26688
rect 18396 26624 18412 26688
rect 18476 26624 18492 26688
rect 18556 26624 18564 26688
rect 18244 25600 18564 26624
rect 18244 25536 18252 25600
rect 18316 25546 18332 25600
rect 18396 25546 18412 25600
rect 18476 25546 18492 25600
rect 18556 25536 18564 25600
rect 18244 25310 18286 25536
rect 18522 25310 18564 25536
rect 18244 24512 18564 25310
rect 18244 24448 18252 24512
rect 18316 24448 18332 24512
rect 18396 24448 18412 24512
rect 18476 24448 18492 24512
rect 18556 24448 18564 24512
rect 18244 23424 18564 24448
rect 18244 23360 18252 23424
rect 18316 23360 18332 23424
rect 18396 23360 18412 23424
rect 18476 23360 18492 23424
rect 18556 23360 18564 23424
rect 18244 22546 18564 23360
rect 18244 22336 18286 22546
rect 18522 22336 18564 22546
rect 18244 22272 18252 22336
rect 18316 22272 18332 22310
rect 18396 22272 18412 22310
rect 18476 22272 18492 22310
rect 18556 22272 18564 22336
rect 18244 21248 18564 22272
rect 18244 21184 18252 21248
rect 18316 21184 18332 21248
rect 18396 21184 18412 21248
rect 18476 21184 18492 21248
rect 18556 21184 18564 21248
rect 18244 20160 18564 21184
rect 18244 20096 18252 20160
rect 18316 20096 18332 20160
rect 18396 20096 18412 20160
rect 18476 20096 18492 20160
rect 18556 20096 18564 20160
rect 18244 19546 18564 20096
rect 18244 19310 18286 19546
rect 18522 19310 18564 19546
rect 18244 19072 18564 19310
rect 18244 19008 18252 19072
rect 18316 19008 18332 19072
rect 18396 19008 18412 19072
rect 18476 19008 18492 19072
rect 18556 19008 18564 19072
rect 18244 17984 18564 19008
rect 18244 17920 18252 17984
rect 18316 17920 18332 17984
rect 18396 17920 18412 17984
rect 18476 17920 18492 17984
rect 18556 17920 18564 17984
rect 18244 16896 18564 17920
rect 18244 16832 18252 16896
rect 18316 16832 18332 16896
rect 18396 16832 18412 16896
rect 18476 16832 18492 16896
rect 18556 16832 18564 16896
rect 18244 16546 18564 16832
rect 18244 16310 18286 16546
rect 18522 16310 18564 16546
rect 18244 15808 18564 16310
rect 18244 15744 18252 15808
rect 18316 15744 18332 15808
rect 18396 15744 18412 15808
rect 18476 15744 18492 15808
rect 18556 15744 18564 15808
rect 18244 14720 18564 15744
rect 18244 14656 18252 14720
rect 18316 14656 18332 14720
rect 18396 14656 18412 14720
rect 18476 14656 18492 14720
rect 18556 14656 18564 14720
rect 18244 13632 18564 14656
rect 18244 13568 18252 13632
rect 18316 13568 18332 13632
rect 18396 13568 18412 13632
rect 18476 13568 18492 13632
rect 18556 13568 18564 13632
rect 18244 13546 18564 13568
rect 18244 13310 18286 13546
rect 18522 13310 18564 13546
rect 18244 12544 18564 13310
rect 18244 12480 18252 12544
rect 18316 12480 18332 12544
rect 18396 12480 18412 12544
rect 18476 12480 18492 12544
rect 18556 12480 18564 12544
rect 18244 11456 18564 12480
rect 18244 11392 18252 11456
rect 18316 11392 18332 11456
rect 18396 11392 18412 11456
rect 18476 11392 18492 11456
rect 18556 11392 18564 11456
rect 18244 10546 18564 11392
rect 18244 10368 18286 10546
rect 18522 10368 18564 10546
rect 18244 10304 18252 10368
rect 18316 10304 18332 10310
rect 18396 10304 18412 10310
rect 18476 10304 18492 10310
rect 18556 10304 18564 10368
rect 18244 9280 18564 10304
rect 18244 9216 18252 9280
rect 18316 9216 18332 9280
rect 18396 9216 18412 9280
rect 18476 9216 18492 9280
rect 18556 9216 18564 9280
rect 18244 8192 18564 9216
rect 18244 8128 18252 8192
rect 18316 8128 18332 8192
rect 18396 8128 18412 8192
rect 18476 8128 18492 8192
rect 18556 8128 18564 8192
rect 18244 7546 18564 8128
rect 18244 7310 18286 7546
rect 18522 7310 18564 7546
rect 18244 7104 18564 7310
rect 18244 7040 18252 7104
rect 18316 7040 18332 7104
rect 18396 7040 18412 7104
rect 18476 7040 18492 7104
rect 18556 7040 18564 7104
rect 18244 6016 18564 7040
rect 18244 5952 18252 6016
rect 18316 5952 18332 6016
rect 18396 5952 18412 6016
rect 18476 5952 18492 6016
rect 18556 5952 18564 6016
rect 18244 4928 18564 5952
rect 18244 4864 18252 4928
rect 18316 4864 18332 4928
rect 18396 4864 18412 4928
rect 18476 4864 18492 4928
rect 18556 4864 18564 4928
rect 18244 4546 18564 4864
rect 18244 4310 18286 4546
rect 18522 4310 18564 4546
rect 18244 3840 18564 4310
rect 18244 3776 18252 3840
rect 18316 3776 18332 3840
rect 18396 3776 18412 3840
rect 18476 3776 18492 3840
rect 18556 3776 18564 3840
rect 18244 2752 18564 3776
rect 18244 2688 18252 2752
rect 18316 2688 18332 2752
rect 18396 2688 18412 2752
rect 18476 2688 18492 2752
rect 18556 2688 18564 2752
rect 18244 2128 18564 2688
rect 19744 29408 20064 29424
rect 19744 29344 19752 29408
rect 19816 29344 19832 29408
rect 19896 29344 19912 29408
rect 19976 29344 19992 29408
rect 20056 29344 20064 29408
rect 19744 28320 20064 29344
rect 19744 28256 19752 28320
rect 19816 28256 19832 28320
rect 19896 28256 19912 28320
rect 19976 28256 19992 28320
rect 20056 28256 20064 28320
rect 19744 27232 20064 28256
rect 19744 27168 19752 27232
rect 19816 27168 19832 27232
rect 19896 27168 19912 27232
rect 19976 27168 19992 27232
rect 20056 27168 20064 27232
rect 19744 27046 20064 27168
rect 19744 26810 19786 27046
rect 20022 26810 20064 27046
rect 19744 26144 20064 26810
rect 19744 26080 19752 26144
rect 19816 26080 19832 26144
rect 19896 26080 19912 26144
rect 19976 26080 19992 26144
rect 20056 26080 20064 26144
rect 19744 25056 20064 26080
rect 19744 24992 19752 25056
rect 19816 24992 19832 25056
rect 19896 24992 19912 25056
rect 19976 24992 19992 25056
rect 20056 24992 20064 25056
rect 19744 24046 20064 24992
rect 19744 23968 19786 24046
rect 20022 23968 20064 24046
rect 19744 23904 19752 23968
rect 20056 23904 20064 23968
rect 19744 23810 19786 23904
rect 20022 23810 20064 23904
rect 19744 22880 20064 23810
rect 19744 22816 19752 22880
rect 19816 22816 19832 22880
rect 19896 22816 19912 22880
rect 19976 22816 19992 22880
rect 20056 22816 20064 22880
rect 19744 21792 20064 22816
rect 19744 21728 19752 21792
rect 19816 21728 19832 21792
rect 19896 21728 19912 21792
rect 19976 21728 19992 21792
rect 20056 21728 20064 21792
rect 19744 21046 20064 21728
rect 19744 20810 19786 21046
rect 20022 20810 20064 21046
rect 19744 20704 20064 20810
rect 19744 20640 19752 20704
rect 19816 20640 19832 20704
rect 19896 20640 19912 20704
rect 19976 20640 19992 20704
rect 20056 20640 20064 20704
rect 19744 19616 20064 20640
rect 19744 19552 19752 19616
rect 19816 19552 19832 19616
rect 19896 19552 19912 19616
rect 19976 19552 19992 19616
rect 20056 19552 20064 19616
rect 19744 18528 20064 19552
rect 19744 18464 19752 18528
rect 19816 18464 19832 18528
rect 19896 18464 19912 18528
rect 19976 18464 19992 18528
rect 20056 18464 20064 18528
rect 19744 18046 20064 18464
rect 19744 17810 19786 18046
rect 20022 17810 20064 18046
rect 19744 17440 20064 17810
rect 19744 17376 19752 17440
rect 19816 17376 19832 17440
rect 19896 17376 19912 17440
rect 19976 17376 19992 17440
rect 20056 17376 20064 17440
rect 19744 16352 20064 17376
rect 19744 16288 19752 16352
rect 19816 16288 19832 16352
rect 19896 16288 19912 16352
rect 19976 16288 19992 16352
rect 20056 16288 20064 16352
rect 19744 15264 20064 16288
rect 19744 15200 19752 15264
rect 19816 15200 19832 15264
rect 19896 15200 19912 15264
rect 19976 15200 19992 15264
rect 20056 15200 20064 15264
rect 19744 15046 20064 15200
rect 19744 14810 19786 15046
rect 20022 14810 20064 15046
rect 19744 14176 20064 14810
rect 19744 14112 19752 14176
rect 19816 14112 19832 14176
rect 19896 14112 19912 14176
rect 19976 14112 19992 14176
rect 20056 14112 20064 14176
rect 19744 13088 20064 14112
rect 19744 13024 19752 13088
rect 19816 13024 19832 13088
rect 19896 13024 19912 13088
rect 19976 13024 19992 13088
rect 20056 13024 20064 13088
rect 19744 12046 20064 13024
rect 19744 12000 19786 12046
rect 20022 12000 20064 12046
rect 19744 11936 19752 12000
rect 20056 11936 20064 12000
rect 19744 11810 19786 11936
rect 20022 11810 20064 11936
rect 19744 10912 20064 11810
rect 19744 10848 19752 10912
rect 19816 10848 19832 10912
rect 19896 10848 19912 10912
rect 19976 10848 19992 10912
rect 20056 10848 20064 10912
rect 19744 9824 20064 10848
rect 19744 9760 19752 9824
rect 19816 9760 19832 9824
rect 19896 9760 19912 9824
rect 19976 9760 19992 9824
rect 20056 9760 20064 9824
rect 19744 9046 20064 9760
rect 19744 8810 19786 9046
rect 20022 8810 20064 9046
rect 19744 8736 20064 8810
rect 19744 8672 19752 8736
rect 19816 8672 19832 8736
rect 19896 8672 19912 8736
rect 19976 8672 19992 8736
rect 20056 8672 20064 8736
rect 19744 7648 20064 8672
rect 19744 7584 19752 7648
rect 19816 7584 19832 7648
rect 19896 7584 19912 7648
rect 19976 7584 19992 7648
rect 20056 7584 20064 7648
rect 19744 6560 20064 7584
rect 19744 6496 19752 6560
rect 19816 6496 19832 6560
rect 19896 6496 19912 6560
rect 19976 6496 19992 6560
rect 20056 6496 20064 6560
rect 19744 6046 20064 6496
rect 19744 5810 19786 6046
rect 20022 5810 20064 6046
rect 19744 5472 20064 5810
rect 19744 5408 19752 5472
rect 19816 5408 19832 5472
rect 19896 5408 19912 5472
rect 19976 5408 19992 5472
rect 20056 5408 20064 5472
rect 19744 4384 20064 5408
rect 19744 4320 19752 4384
rect 19816 4320 19832 4384
rect 19896 4320 19912 4384
rect 19976 4320 19992 4384
rect 20056 4320 20064 4384
rect 19744 3296 20064 4320
rect 19744 3232 19752 3296
rect 19816 3232 19832 3296
rect 19896 3232 19912 3296
rect 19976 3232 19992 3296
rect 20056 3232 20064 3296
rect 19744 3046 20064 3232
rect 19744 2810 19786 3046
rect 20022 2810 20064 3046
rect 19744 2208 20064 2810
rect 19744 2144 19752 2208
rect 19816 2144 19832 2208
rect 19896 2144 19912 2208
rect 19976 2144 19992 2208
rect 20056 2144 20064 2208
rect 19744 2128 20064 2144
rect 21244 28864 21564 29424
rect 21244 28800 21252 28864
rect 21316 28800 21332 28864
rect 21396 28800 21412 28864
rect 21476 28800 21492 28864
rect 21556 28800 21564 28864
rect 21244 28546 21564 28800
rect 21244 28310 21286 28546
rect 21522 28310 21564 28546
rect 21244 27776 21564 28310
rect 21244 27712 21252 27776
rect 21316 27712 21332 27776
rect 21396 27712 21412 27776
rect 21476 27712 21492 27776
rect 21556 27712 21564 27776
rect 21244 26688 21564 27712
rect 21244 26624 21252 26688
rect 21316 26624 21332 26688
rect 21396 26624 21412 26688
rect 21476 26624 21492 26688
rect 21556 26624 21564 26688
rect 21244 25600 21564 26624
rect 21244 25536 21252 25600
rect 21316 25546 21332 25600
rect 21396 25546 21412 25600
rect 21476 25546 21492 25600
rect 21556 25536 21564 25600
rect 21244 25310 21286 25536
rect 21522 25310 21564 25536
rect 21244 24512 21564 25310
rect 21244 24448 21252 24512
rect 21316 24448 21332 24512
rect 21396 24448 21412 24512
rect 21476 24448 21492 24512
rect 21556 24448 21564 24512
rect 21244 23424 21564 24448
rect 21244 23360 21252 23424
rect 21316 23360 21332 23424
rect 21396 23360 21412 23424
rect 21476 23360 21492 23424
rect 21556 23360 21564 23424
rect 21244 22546 21564 23360
rect 21244 22336 21286 22546
rect 21522 22336 21564 22546
rect 21244 22272 21252 22336
rect 21316 22272 21332 22310
rect 21396 22272 21412 22310
rect 21476 22272 21492 22310
rect 21556 22272 21564 22336
rect 21244 21248 21564 22272
rect 21244 21184 21252 21248
rect 21316 21184 21332 21248
rect 21396 21184 21412 21248
rect 21476 21184 21492 21248
rect 21556 21184 21564 21248
rect 21244 20160 21564 21184
rect 21244 20096 21252 20160
rect 21316 20096 21332 20160
rect 21396 20096 21412 20160
rect 21476 20096 21492 20160
rect 21556 20096 21564 20160
rect 21244 19546 21564 20096
rect 21244 19310 21286 19546
rect 21522 19310 21564 19546
rect 21244 19072 21564 19310
rect 21244 19008 21252 19072
rect 21316 19008 21332 19072
rect 21396 19008 21412 19072
rect 21476 19008 21492 19072
rect 21556 19008 21564 19072
rect 21244 17984 21564 19008
rect 21244 17920 21252 17984
rect 21316 17920 21332 17984
rect 21396 17920 21412 17984
rect 21476 17920 21492 17984
rect 21556 17920 21564 17984
rect 21244 16896 21564 17920
rect 21244 16832 21252 16896
rect 21316 16832 21332 16896
rect 21396 16832 21412 16896
rect 21476 16832 21492 16896
rect 21556 16832 21564 16896
rect 21244 16546 21564 16832
rect 21244 16310 21286 16546
rect 21522 16310 21564 16546
rect 21244 15808 21564 16310
rect 21244 15744 21252 15808
rect 21316 15744 21332 15808
rect 21396 15744 21412 15808
rect 21476 15744 21492 15808
rect 21556 15744 21564 15808
rect 21244 14720 21564 15744
rect 21244 14656 21252 14720
rect 21316 14656 21332 14720
rect 21396 14656 21412 14720
rect 21476 14656 21492 14720
rect 21556 14656 21564 14720
rect 21244 13632 21564 14656
rect 21244 13568 21252 13632
rect 21316 13568 21332 13632
rect 21396 13568 21412 13632
rect 21476 13568 21492 13632
rect 21556 13568 21564 13632
rect 21244 13546 21564 13568
rect 21244 13310 21286 13546
rect 21522 13310 21564 13546
rect 21244 12544 21564 13310
rect 21244 12480 21252 12544
rect 21316 12480 21332 12544
rect 21396 12480 21412 12544
rect 21476 12480 21492 12544
rect 21556 12480 21564 12544
rect 21244 11456 21564 12480
rect 21244 11392 21252 11456
rect 21316 11392 21332 11456
rect 21396 11392 21412 11456
rect 21476 11392 21492 11456
rect 21556 11392 21564 11456
rect 21244 10546 21564 11392
rect 21244 10368 21286 10546
rect 21522 10368 21564 10546
rect 21244 10304 21252 10368
rect 21316 10304 21332 10310
rect 21396 10304 21412 10310
rect 21476 10304 21492 10310
rect 21556 10304 21564 10368
rect 21244 9280 21564 10304
rect 21244 9216 21252 9280
rect 21316 9216 21332 9280
rect 21396 9216 21412 9280
rect 21476 9216 21492 9280
rect 21556 9216 21564 9280
rect 21244 8192 21564 9216
rect 21244 8128 21252 8192
rect 21316 8128 21332 8192
rect 21396 8128 21412 8192
rect 21476 8128 21492 8192
rect 21556 8128 21564 8192
rect 21244 7546 21564 8128
rect 21244 7310 21286 7546
rect 21522 7310 21564 7546
rect 21244 7104 21564 7310
rect 21244 7040 21252 7104
rect 21316 7040 21332 7104
rect 21396 7040 21412 7104
rect 21476 7040 21492 7104
rect 21556 7040 21564 7104
rect 21244 6016 21564 7040
rect 21244 5952 21252 6016
rect 21316 5952 21332 6016
rect 21396 5952 21412 6016
rect 21476 5952 21492 6016
rect 21556 5952 21564 6016
rect 21244 4928 21564 5952
rect 21244 4864 21252 4928
rect 21316 4864 21332 4928
rect 21396 4864 21412 4928
rect 21476 4864 21492 4928
rect 21556 4864 21564 4928
rect 21244 4546 21564 4864
rect 21244 4310 21286 4546
rect 21522 4310 21564 4546
rect 21244 3840 21564 4310
rect 21244 3776 21252 3840
rect 21316 3776 21332 3840
rect 21396 3776 21412 3840
rect 21476 3776 21492 3840
rect 21556 3776 21564 3840
rect 21244 2752 21564 3776
rect 21244 2688 21252 2752
rect 21316 2688 21332 2752
rect 21396 2688 21412 2752
rect 21476 2688 21492 2752
rect 21556 2688 21564 2752
rect 21244 2128 21564 2688
rect 22744 29408 23064 29424
rect 22744 29344 22752 29408
rect 22816 29344 22832 29408
rect 22896 29344 22912 29408
rect 22976 29344 22992 29408
rect 23056 29344 23064 29408
rect 22744 28320 23064 29344
rect 22744 28256 22752 28320
rect 22816 28256 22832 28320
rect 22896 28256 22912 28320
rect 22976 28256 22992 28320
rect 23056 28256 23064 28320
rect 22744 27232 23064 28256
rect 22744 27168 22752 27232
rect 22816 27168 22832 27232
rect 22896 27168 22912 27232
rect 22976 27168 22992 27232
rect 23056 27168 23064 27232
rect 22744 27046 23064 27168
rect 22744 26810 22786 27046
rect 23022 26810 23064 27046
rect 22744 26144 23064 26810
rect 22744 26080 22752 26144
rect 22816 26080 22832 26144
rect 22896 26080 22912 26144
rect 22976 26080 22992 26144
rect 23056 26080 23064 26144
rect 22744 25056 23064 26080
rect 22744 24992 22752 25056
rect 22816 24992 22832 25056
rect 22896 24992 22912 25056
rect 22976 24992 22992 25056
rect 23056 24992 23064 25056
rect 22744 24046 23064 24992
rect 22744 23968 22786 24046
rect 23022 23968 23064 24046
rect 22744 23904 22752 23968
rect 23056 23904 23064 23968
rect 22744 23810 22786 23904
rect 23022 23810 23064 23904
rect 22744 22880 23064 23810
rect 22744 22816 22752 22880
rect 22816 22816 22832 22880
rect 22896 22816 22912 22880
rect 22976 22816 22992 22880
rect 23056 22816 23064 22880
rect 22744 21792 23064 22816
rect 22744 21728 22752 21792
rect 22816 21728 22832 21792
rect 22896 21728 22912 21792
rect 22976 21728 22992 21792
rect 23056 21728 23064 21792
rect 22744 21046 23064 21728
rect 22744 20810 22786 21046
rect 23022 20810 23064 21046
rect 22744 20704 23064 20810
rect 22744 20640 22752 20704
rect 22816 20640 22832 20704
rect 22896 20640 22912 20704
rect 22976 20640 22992 20704
rect 23056 20640 23064 20704
rect 22744 19616 23064 20640
rect 22744 19552 22752 19616
rect 22816 19552 22832 19616
rect 22896 19552 22912 19616
rect 22976 19552 22992 19616
rect 23056 19552 23064 19616
rect 22744 18528 23064 19552
rect 22744 18464 22752 18528
rect 22816 18464 22832 18528
rect 22896 18464 22912 18528
rect 22976 18464 22992 18528
rect 23056 18464 23064 18528
rect 22744 18046 23064 18464
rect 22744 17810 22786 18046
rect 23022 17810 23064 18046
rect 22744 17440 23064 17810
rect 22744 17376 22752 17440
rect 22816 17376 22832 17440
rect 22896 17376 22912 17440
rect 22976 17376 22992 17440
rect 23056 17376 23064 17440
rect 22744 16352 23064 17376
rect 22744 16288 22752 16352
rect 22816 16288 22832 16352
rect 22896 16288 22912 16352
rect 22976 16288 22992 16352
rect 23056 16288 23064 16352
rect 22744 15264 23064 16288
rect 22744 15200 22752 15264
rect 22816 15200 22832 15264
rect 22896 15200 22912 15264
rect 22976 15200 22992 15264
rect 23056 15200 23064 15264
rect 22744 15046 23064 15200
rect 22744 14810 22786 15046
rect 23022 14810 23064 15046
rect 22744 14176 23064 14810
rect 22744 14112 22752 14176
rect 22816 14112 22832 14176
rect 22896 14112 22912 14176
rect 22976 14112 22992 14176
rect 23056 14112 23064 14176
rect 22744 13088 23064 14112
rect 22744 13024 22752 13088
rect 22816 13024 22832 13088
rect 22896 13024 22912 13088
rect 22976 13024 22992 13088
rect 23056 13024 23064 13088
rect 22744 12046 23064 13024
rect 22744 12000 22786 12046
rect 23022 12000 23064 12046
rect 22744 11936 22752 12000
rect 23056 11936 23064 12000
rect 22744 11810 22786 11936
rect 23022 11810 23064 11936
rect 22744 10912 23064 11810
rect 22744 10848 22752 10912
rect 22816 10848 22832 10912
rect 22896 10848 22912 10912
rect 22976 10848 22992 10912
rect 23056 10848 23064 10912
rect 22744 9824 23064 10848
rect 22744 9760 22752 9824
rect 22816 9760 22832 9824
rect 22896 9760 22912 9824
rect 22976 9760 22992 9824
rect 23056 9760 23064 9824
rect 22744 9046 23064 9760
rect 22744 8810 22786 9046
rect 23022 8810 23064 9046
rect 22744 8736 23064 8810
rect 22744 8672 22752 8736
rect 22816 8672 22832 8736
rect 22896 8672 22912 8736
rect 22976 8672 22992 8736
rect 23056 8672 23064 8736
rect 22744 7648 23064 8672
rect 22744 7584 22752 7648
rect 22816 7584 22832 7648
rect 22896 7584 22912 7648
rect 22976 7584 22992 7648
rect 23056 7584 23064 7648
rect 22744 6560 23064 7584
rect 22744 6496 22752 6560
rect 22816 6496 22832 6560
rect 22896 6496 22912 6560
rect 22976 6496 22992 6560
rect 23056 6496 23064 6560
rect 22744 6046 23064 6496
rect 22744 5810 22786 6046
rect 23022 5810 23064 6046
rect 22744 5472 23064 5810
rect 22744 5408 22752 5472
rect 22816 5408 22832 5472
rect 22896 5408 22912 5472
rect 22976 5408 22992 5472
rect 23056 5408 23064 5472
rect 22744 4384 23064 5408
rect 22744 4320 22752 4384
rect 22816 4320 22832 4384
rect 22896 4320 22912 4384
rect 22976 4320 22992 4384
rect 23056 4320 23064 4384
rect 22744 3296 23064 4320
rect 22744 3232 22752 3296
rect 22816 3232 22832 3296
rect 22896 3232 22912 3296
rect 22976 3232 22992 3296
rect 23056 3232 23064 3296
rect 22744 3046 23064 3232
rect 22744 2810 22786 3046
rect 23022 2810 23064 3046
rect 22744 2208 23064 2810
rect 22744 2144 22752 2208
rect 22816 2144 22832 2208
rect 22896 2144 22912 2208
rect 22976 2144 22992 2208
rect 23056 2144 23064 2208
rect 22744 2128 23064 2144
rect 24244 28864 24564 29424
rect 24244 28800 24252 28864
rect 24316 28800 24332 28864
rect 24396 28800 24412 28864
rect 24476 28800 24492 28864
rect 24556 28800 24564 28864
rect 24244 28546 24564 28800
rect 24244 28310 24286 28546
rect 24522 28310 24564 28546
rect 24244 27776 24564 28310
rect 24244 27712 24252 27776
rect 24316 27712 24332 27776
rect 24396 27712 24412 27776
rect 24476 27712 24492 27776
rect 24556 27712 24564 27776
rect 24244 26688 24564 27712
rect 24244 26624 24252 26688
rect 24316 26624 24332 26688
rect 24396 26624 24412 26688
rect 24476 26624 24492 26688
rect 24556 26624 24564 26688
rect 24244 25600 24564 26624
rect 24244 25536 24252 25600
rect 24316 25546 24332 25600
rect 24396 25546 24412 25600
rect 24476 25546 24492 25600
rect 24556 25536 24564 25600
rect 24244 25310 24286 25536
rect 24522 25310 24564 25536
rect 24244 24512 24564 25310
rect 24244 24448 24252 24512
rect 24316 24448 24332 24512
rect 24396 24448 24412 24512
rect 24476 24448 24492 24512
rect 24556 24448 24564 24512
rect 24244 23424 24564 24448
rect 24244 23360 24252 23424
rect 24316 23360 24332 23424
rect 24396 23360 24412 23424
rect 24476 23360 24492 23424
rect 24556 23360 24564 23424
rect 24244 22546 24564 23360
rect 24244 22336 24286 22546
rect 24522 22336 24564 22546
rect 24244 22272 24252 22336
rect 24316 22272 24332 22310
rect 24396 22272 24412 22310
rect 24476 22272 24492 22310
rect 24556 22272 24564 22336
rect 24244 21248 24564 22272
rect 24244 21184 24252 21248
rect 24316 21184 24332 21248
rect 24396 21184 24412 21248
rect 24476 21184 24492 21248
rect 24556 21184 24564 21248
rect 24244 20160 24564 21184
rect 24244 20096 24252 20160
rect 24316 20096 24332 20160
rect 24396 20096 24412 20160
rect 24476 20096 24492 20160
rect 24556 20096 24564 20160
rect 24244 19546 24564 20096
rect 24244 19310 24286 19546
rect 24522 19310 24564 19546
rect 24244 19072 24564 19310
rect 24244 19008 24252 19072
rect 24316 19008 24332 19072
rect 24396 19008 24412 19072
rect 24476 19008 24492 19072
rect 24556 19008 24564 19072
rect 24244 17984 24564 19008
rect 24244 17920 24252 17984
rect 24316 17920 24332 17984
rect 24396 17920 24412 17984
rect 24476 17920 24492 17984
rect 24556 17920 24564 17984
rect 24244 16896 24564 17920
rect 24244 16832 24252 16896
rect 24316 16832 24332 16896
rect 24396 16832 24412 16896
rect 24476 16832 24492 16896
rect 24556 16832 24564 16896
rect 24244 16546 24564 16832
rect 24244 16310 24286 16546
rect 24522 16310 24564 16546
rect 24244 15808 24564 16310
rect 24244 15744 24252 15808
rect 24316 15744 24332 15808
rect 24396 15744 24412 15808
rect 24476 15744 24492 15808
rect 24556 15744 24564 15808
rect 24244 14720 24564 15744
rect 24244 14656 24252 14720
rect 24316 14656 24332 14720
rect 24396 14656 24412 14720
rect 24476 14656 24492 14720
rect 24556 14656 24564 14720
rect 24244 13632 24564 14656
rect 24244 13568 24252 13632
rect 24316 13568 24332 13632
rect 24396 13568 24412 13632
rect 24476 13568 24492 13632
rect 24556 13568 24564 13632
rect 24244 13546 24564 13568
rect 24244 13310 24286 13546
rect 24522 13310 24564 13546
rect 24244 12544 24564 13310
rect 24244 12480 24252 12544
rect 24316 12480 24332 12544
rect 24396 12480 24412 12544
rect 24476 12480 24492 12544
rect 24556 12480 24564 12544
rect 24244 11456 24564 12480
rect 24244 11392 24252 11456
rect 24316 11392 24332 11456
rect 24396 11392 24412 11456
rect 24476 11392 24492 11456
rect 24556 11392 24564 11456
rect 24244 10546 24564 11392
rect 24244 10368 24286 10546
rect 24522 10368 24564 10546
rect 24244 10304 24252 10368
rect 24316 10304 24332 10310
rect 24396 10304 24412 10310
rect 24476 10304 24492 10310
rect 24556 10304 24564 10368
rect 24244 9280 24564 10304
rect 24244 9216 24252 9280
rect 24316 9216 24332 9280
rect 24396 9216 24412 9280
rect 24476 9216 24492 9280
rect 24556 9216 24564 9280
rect 24244 8192 24564 9216
rect 24244 8128 24252 8192
rect 24316 8128 24332 8192
rect 24396 8128 24412 8192
rect 24476 8128 24492 8192
rect 24556 8128 24564 8192
rect 24244 7546 24564 8128
rect 24244 7310 24286 7546
rect 24522 7310 24564 7546
rect 24244 7104 24564 7310
rect 24244 7040 24252 7104
rect 24316 7040 24332 7104
rect 24396 7040 24412 7104
rect 24476 7040 24492 7104
rect 24556 7040 24564 7104
rect 24244 6016 24564 7040
rect 24244 5952 24252 6016
rect 24316 5952 24332 6016
rect 24396 5952 24412 6016
rect 24476 5952 24492 6016
rect 24556 5952 24564 6016
rect 24244 4928 24564 5952
rect 24244 4864 24252 4928
rect 24316 4864 24332 4928
rect 24396 4864 24412 4928
rect 24476 4864 24492 4928
rect 24556 4864 24564 4928
rect 24244 4546 24564 4864
rect 24244 4310 24286 4546
rect 24522 4310 24564 4546
rect 24244 3840 24564 4310
rect 24244 3776 24252 3840
rect 24316 3776 24332 3840
rect 24396 3776 24412 3840
rect 24476 3776 24492 3840
rect 24556 3776 24564 3840
rect 24244 2752 24564 3776
rect 24244 2688 24252 2752
rect 24316 2688 24332 2752
rect 24396 2688 24412 2752
rect 24476 2688 24492 2752
rect 24556 2688 24564 2752
rect 24244 2128 24564 2688
rect 25744 29408 26064 29424
rect 25744 29344 25752 29408
rect 25816 29344 25832 29408
rect 25896 29344 25912 29408
rect 25976 29344 25992 29408
rect 26056 29344 26064 29408
rect 25744 28320 26064 29344
rect 25744 28256 25752 28320
rect 25816 28256 25832 28320
rect 25896 28256 25912 28320
rect 25976 28256 25992 28320
rect 26056 28256 26064 28320
rect 25744 27232 26064 28256
rect 25744 27168 25752 27232
rect 25816 27168 25832 27232
rect 25896 27168 25912 27232
rect 25976 27168 25992 27232
rect 26056 27168 26064 27232
rect 25744 27046 26064 27168
rect 25744 26810 25786 27046
rect 26022 26810 26064 27046
rect 25744 26144 26064 26810
rect 25744 26080 25752 26144
rect 25816 26080 25832 26144
rect 25896 26080 25912 26144
rect 25976 26080 25992 26144
rect 26056 26080 26064 26144
rect 25744 25056 26064 26080
rect 25744 24992 25752 25056
rect 25816 24992 25832 25056
rect 25896 24992 25912 25056
rect 25976 24992 25992 25056
rect 26056 24992 26064 25056
rect 25744 24046 26064 24992
rect 25744 23968 25786 24046
rect 26022 23968 26064 24046
rect 25744 23904 25752 23968
rect 26056 23904 26064 23968
rect 25744 23810 25786 23904
rect 26022 23810 26064 23904
rect 25744 22880 26064 23810
rect 25744 22816 25752 22880
rect 25816 22816 25832 22880
rect 25896 22816 25912 22880
rect 25976 22816 25992 22880
rect 26056 22816 26064 22880
rect 25744 21792 26064 22816
rect 25744 21728 25752 21792
rect 25816 21728 25832 21792
rect 25896 21728 25912 21792
rect 25976 21728 25992 21792
rect 26056 21728 26064 21792
rect 25744 21046 26064 21728
rect 25744 20810 25786 21046
rect 26022 20810 26064 21046
rect 25744 20704 26064 20810
rect 25744 20640 25752 20704
rect 25816 20640 25832 20704
rect 25896 20640 25912 20704
rect 25976 20640 25992 20704
rect 26056 20640 26064 20704
rect 25744 19616 26064 20640
rect 25744 19552 25752 19616
rect 25816 19552 25832 19616
rect 25896 19552 25912 19616
rect 25976 19552 25992 19616
rect 26056 19552 26064 19616
rect 25744 18528 26064 19552
rect 25744 18464 25752 18528
rect 25816 18464 25832 18528
rect 25896 18464 25912 18528
rect 25976 18464 25992 18528
rect 26056 18464 26064 18528
rect 25744 18046 26064 18464
rect 25744 17810 25786 18046
rect 26022 17810 26064 18046
rect 25744 17440 26064 17810
rect 25744 17376 25752 17440
rect 25816 17376 25832 17440
rect 25896 17376 25912 17440
rect 25976 17376 25992 17440
rect 26056 17376 26064 17440
rect 25744 16352 26064 17376
rect 25744 16288 25752 16352
rect 25816 16288 25832 16352
rect 25896 16288 25912 16352
rect 25976 16288 25992 16352
rect 26056 16288 26064 16352
rect 25744 15264 26064 16288
rect 25744 15200 25752 15264
rect 25816 15200 25832 15264
rect 25896 15200 25912 15264
rect 25976 15200 25992 15264
rect 26056 15200 26064 15264
rect 25744 15046 26064 15200
rect 25744 14810 25786 15046
rect 26022 14810 26064 15046
rect 25744 14176 26064 14810
rect 25744 14112 25752 14176
rect 25816 14112 25832 14176
rect 25896 14112 25912 14176
rect 25976 14112 25992 14176
rect 26056 14112 26064 14176
rect 25744 13088 26064 14112
rect 25744 13024 25752 13088
rect 25816 13024 25832 13088
rect 25896 13024 25912 13088
rect 25976 13024 25992 13088
rect 26056 13024 26064 13088
rect 25744 12046 26064 13024
rect 25744 12000 25786 12046
rect 26022 12000 26064 12046
rect 25744 11936 25752 12000
rect 26056 11936 26064 12000
rect 25744 11810 25786 11936
rect 26022 11810 26064 11936
rect 25744 10912 26064 11810
rect 25744 10848 25752 10912
rect 25816 10848 25832 10912
rect 25896 10848 25912 10912
rect 25976 10848 25992 10912
rect 26056 10848 26064 10912
rect 25744 9824 26064 10848
rect 25744 9760 25752 9824
rect 25816 9760 25832 9824
rect 25896 9760 25912 9824
rect 25976 9760 25992 9824
rect 26056 9760 26064 9824
rect 25744 9046 26064 9760
rect 25744 8810 25786 9046
rect 26022 8810 26064 9046
rect 25744 8736 26064 8810
rect 25744 8672 25752 8736
rect 25816 8672 25832 8736
rect 25896 8672 25912 8736
rect 25976 8672 25992 8736
rect 26056 8672 26064 8736
rect 25744 7648 26064 8672
rect 25744 7584 25752 7648
rect 25816 7584 25832 7648
rect 25896 7584 25912 7648
rect 25976 7584 25992 7648
rect 26056 7584 26064 7648
rect 25744 6560 26064 7584
rect 25744 6496 25752 6560
rect 25816 6496 25832 6560
rect 25896 6496 25912 6560
rect 25976 6496 25992 6560
rect 26056 6496 26064 6560
rect 25744 6046 26064 6496
rect 25744 5810 25786 6046
rect 26022 5810 26064 6046
rect 25744 5472 26064 5810
rect 25744 5408 25752 5472
rect 25816 5408 25832 5472
rect 25896 5408 25912 5472
rect 25976 5408 25992 5472
rect 26056 5408 26064 5472
rect 25744 4384 26064 5408
rect 25744 4320 25752 4384
rect 25816 4320 25832 4384
rect 25896 4320 25912 4384
rect 25976 4320 25992 4384
rect 26056 4320 26064 4384
rect 25744 3296 26064 4320
rect 25744 3232 25752 3296
rect 25816 3232 25832 3296
rect 25896 3232 25912 3296
rect 25976 3232 25992 3296
rect 26056 3232 26064 3296
rect 25744 3046 26064 3232
rect 25744 2810 25786 3046
rect 26022 2810 26064 3046
rect 25744 2208 26064 2810
rect 25744 2144 25752 2208
rect 25816 2144 25832 2208
rect 25896 2144 25912 2208
rect 25976 2144 25992 2208
rect 26056 2144 26064 2208
rect 25744 2128 26064 2144
rect 27244 28864 27564 29424
rect 27244 28800 27252 28864
rect 27316 28800 27332 28864
rect 27396 28800 27412 28864
rect 27476 28800 27492 28864
rect 27556 28800 27564 28864
rect 27244 28546 27564 28800
rect 27244 28310 27286 28546
rect 27522 28310 27564 28546
rect 27244 27776 27564 28310
rect 27244 27712 27252 27776
rect 27316 27712 27332 27776
rect 27396 27712 27412 27776
rect 27476 27712 27492 27776
rect 27556 27712 27564 27776
rect 27244 26688 27564 27712
rect 27244 26624 27252 26688
rect 27316 26624 27332 26688
rect 27396 26624 27412 26688
rect 27476 26624 27492 26688
rect 27556 26624 27564 26688
rect 27244 25600 27564 26624
rect 27244 25536 27252 25600
rect 27316 25546 27332 25600
rect 27396 25546 27412 25600
rect 27476 25546 27492 25600
rect 27556 25536 27564 25600
rect 27244 25310 27286 25536
rect 27522 25310 27564 25536
rect 27244 24512 27564 25310
rect 27244 24448 27252 24512
rect 27316 24448 27332 24512
rect 27396 24448 27412 24512
rect 27476 24448 27492 24512
rect 27556 24448 27564 24512
rect 27244 23424 27564 24448
rect 27244 23360 27252 23424
rect 27316 23360 27332 23424
rect 27396 23360 27412 23424
rect 27476 23360 27492 23424
rect 27556 23360 27564 23424
rect 27244 22546 27564 23360
rect 27244 22336 27286 22546
rect 27522 22336 27564 22546
rect 27244 22272 27252 22336
rect 27316 22272 27332 22310
rect 27396 22272 27412 22310
rect 27476 22272 27492 22310
rect 27556 22272 27564 22336
rect 27244 21248 27564 22272
rect 27244 21184 27252 21248
rect 27316 21184 27332 21248
rect 27396 21184 27412 21248
rect 27476 21184 27492 21248
rect 27556 21184 27564 21248
rect 27244 20160 27564 21184
rect 27244 20096 27252 20160
rect 27316 20096 27332 20160
rect 27396 20096 27412 20160
rect 27476 20096 27492 20160
rect 27556 20096 27564 20160
rect 27244 19546 27564 20096
rect 27244 19310 27286 19546
rect 27522 19310 27564 19546
rect 27244 19072 27564 19310
rect 27244 19008 27252 19072
rect 27316 19008 27332 19072
rect 27396 19008 27412 19072
rect 27476 19008 27492 19072
rect 27556 19008 27564 19072
rect 27244 17984 27564 19008
rect 27244 17920 27252 17984
rect 27316 17920 27332 17984
rect 27396 17920 27412 17984
rect 27476 17920 27492 17984
rect 27556 17920 27564 17984
rect 27244 16896 27564 17920
rect 27244 16832 27252 16896
rect 27316 16832 27332 16896
rect 27396 16832 27412 16896
rect 27476 16832 27492 16896
rect 27556 16832 27564 16896
rect 27244 16546 27564 16832
rect 27244 16310 27286 16546
rect 27522 16310 27564 16546
rect 27244 15808 27564 16310
rect 27244 15744 27252 15808
rect 27316 15744 27332 15808
rect 27396 15744 27412 15808
rect 27476 15744 27492 15808
rect 27556 15744 27564 15808
rect 27244 14720 27564 15744
rect 27244 14656 27252 14720
rect 27316 14656 27332 14720
rect 27396 14656 27412 14720
rect 27476 14656 27492 14720
rect 27556 14656 27564 14720
rect 27244 13632 27564 14656
rect 27244 13568 27252 13632
rect 27316 13568 27332 13632
rect 27396 13568 27412 13632
rect 27476 13568 27492 13632
rect 27556 13568 27564 13632
rect 27244 13546 27564 13568
rect 27244 13310 27286 13546
rect 27522 13310 27564 13546
rect 27244 12544 27564 13310
rect 27244 12480 27252 12544
rect 27316 12480 27332 12544
rect 27396 12480 27412 12544
rect 27476 12480 27492 12544
rect 27556 12480 27564 12544
rect 27244 11456 27564 12480
rect 27244 11392 27252 11456
rect 27316 11392 27332 11456
rect 27396 11392 27412 11456
rect 27476 11392 27492 11456
rect 27556 11392 27564 11456
rect 27244 10546 27564 11392
rect 27244 10368 27286 10546
rect 27522 10368 27564 10546
rect 27244 10304 27252 10368
rect 27316 10304 27332 10310
rect 27396 10304 27412 10310
rect 27476 10304 27492 10310
rect 27556 10304 27564 10368
rect 27244 9280 27564 10304
rect 27244 9216 27252 9280
rect 27316 9216 27332 9280
rect 27396 9216 27412 9280
rect 27476 9216 27492 9280
rect 27556 9216 27564 9280
rect 27244 8192 27564 9216
rect 27244 8128 27252 8192
rect 27316 8128 27332 8192
rect 27396 8128 27412 8192
rect 27476 8128 27492 8192
rect 27556 8128 27564 8192
rect 27244 7546 27564 8128
rect 27244 7310 27286 7546
rect 27522 7310 27564 7546
rect 27244 7104 27564 7310
rect 27244 7040 27252 7104
rect 27316 7040 27332 7104
rect 27396 7040 27412 7104
rect 27476 7040 27492 7104
rect 27556 7040 27564 7104
rect 27244 6016 27564 7040
rect 27244 5952 27252 6016
rect 27316 5952 27332 6016
rect 27396 5952 27412 6016
rect 27476 5952 27492 6016
rect 27556 5952 27564 6016
rect 27244 4928 27564 5952
rect 27244 4864 27252 4928
rect 27316 4864 27332 4928
rect 27396 4864 27412 4928
rect 27476 4864 27492 4928
rect 27556 4864 27564 4928
rect 27244 4546 27564 4864
rect 27244 4310 27286 4546
rect 27522 4310 27564 4546
rect 27244 3840 27564 4310
rect 27244 3776 27252 3840
rect 27316 3776 27332 3840
rect 27396 3776 27412 3840
rect 27476 3776 27492 3840
rect 27556 3776 27564 3840
rect 27244 2752 27564 3776
rect 27244 2688 27252 2752
rect 27316 2688 27332 2752
rect 27396 2688 27412 2752
rect 27476 2688 27492 2752
rect 27556 2688 27564 2752
rect 27244 2128 27564 2688
<< via4 >>
rect 1786 26810 2022 27046
rect 1786 23968 2022 24046
rect 1786 23904 1816 23968
rect 1816 23904 1832 23968
rect 1832 23904 1896 23968
rect 1896 23904 1912 23968
rect 1912 23904 1976 23968
rect 1976 23904 1992 23968
rect 1992 23904 2022 23968
rect 1786 23810 2022 23904
rect 1786 20810 2022 21046
rect 1786 17810 2022 18046
rect 1786 14810 2022 15046
rect 1786 12000 2022 12046
rect 1786 11936 1816 12000
rect 1816 11936 1832 12000
rect 1832 11936 1896 12000
rect 1896 11936 1912 12000
rect 1912 11936 1976 12000
rect 1976 11936 1992 12000
rect 1992 11936 2022 12000
rect 1786 11810 2022 11936
rect 1786 8810 2022 9046
rect 1786 5810 2022 6046
rect 1786 2810 2022 3046
rect 3286 28310 3522 28546
rect 3286 25536 3316 25546
rect 3316 25536 3332 25546
rect 3332 25536 3396 25546
rect 3396 25536 3412 25546
rect 3412 25536 3476 25546
rect 3476 25536 3492 25546
rect 3492 25536 3522 25546
rect 3286 25310 3522 25536
rect 3286 22336 3522 22546
rect 3286 22310 3316 22336
rect 3316 22310 3332 22336
rect 3332 22310 3396 22336
rect 3396 22310 3412 22336
rect 3412 22310 3476 22336
rect 3476 22310 3492 22336
rect 3492 22310 3522 22336
rect 3286 19310 3522 19546
rect 3286 16310 3522 16546
rect 3286 13310 3522 13546
rect 3286 10368 3522 10546
rect 3286 10310 3316 10368
rect 3316 10310 3332 10368
rect 3332 10310 3396 10368
rect 3396 10310 3412 10368
rect 3412 10310 3476 10368
rect 3476 10310 3492 10368
rect 3492 10310 3522 10368
rect 3286 7310 3522 7546
rect 3286 4310 3522 4546
rect 4786 26810 5022 27046
rect 4786 23968 5022 24046
rect 4786 23904 4816 23968
rect 4816 23904 4832 23968
rect 4832 23904 4896 23968
rect 4896 23904 4912 23968
rect 4912 23904 4976 23968
rect 4976 23904 4992 23968
rect 4992 23904 5022 23968
rect 4786 23810 5022 23904
rect 4786 20810 5022 21046
rect 4786 17810 5022 18046
rect 4786 14810 5022 15046
rect 4786 12000 5022 12046
rect 4786 11936 4816 12000
rect 4816 11936 4832 12000
rect 4832 11936 4896 12000
rect 4896 11936 4912 12000
rect 4912 11936 4976 12000
rect 4976 11936 4992 12000
rect 4992 11936 5022 12000
rect 4786 11810 5022 11936
rect 4786 8810 5022 9046
rect 4786 5810 5022 6046
rect 4786 2810 5022 3046
rect 6286 28310 6522 28546
rect 6286 25536 6316 25546
rect 6316 25536 6332 25546
rect 6332 25536 6396 25546
rect 6396 25536 6412 25546
rect 6412 25536 6476 25546
rect 6476 25536 6492 25546
rect 6492 25536 6522 25546
rect 6286 25310 6522 25536
rect 6286 22336 6522 22546
rect 6286 22310 6316 22336
rect 6316 22310 6332 22336
rect 6332 22310 6396 22336
rect 6396 22310 6412 22336
rect 6412 22310 6476 22336
rect 6476 22310 6492 22336
rect 6492 22310 6522 22336
rect 6286 19310 6522 19546
rect 6286 16310 6522 16546
rect 6286 13310 6522 13546
rect 6286 10368 6522 10546
rect 6286 10310 6316 10368
rect 6316 10310 6332 10368
rect 6332 10310 6396 10368
rect 6396 10310 6412 10368
rect 6412 10310 6476 10368
rect 6476 10310 6492 10368
rect 6492 10310 6522 10368
rect 6286 7310 6522 7546
rect 6286 4310 6522 4546
rect 7786 26810 8022 27046
rect 7786 23968 8022 24046
rect 7786 23904 7816 23968
rect 7816 23904 7832 23968
rect 7832 23904 7896 23968
rect 7896 23904 7912 23968
rect 7912 23904 7976 23968
rect 7976 23904 7992 23968
rect 7992 23904 8022 23968
rect 7786 23810 8022 23904
rect 7786 20810 8022 21046
rect 7786 17810 8022 18046
rect 7786 14810 8022 15046
rect 7786 12000 8022 12046
rect 7786 11936 7816 12000
rect 7816 11936 7832 12000
rect 7832 11936 7896 12000
rect 7896 11936 7912 12000
rect 7912 11936 7976 12000
rect 7976 11936 7992 12000
rect 7992 11936 8022 12000
rect 7786 11810 8022 11936
rect 7786 8810 8022 9046
rect 7786 5810 8022 6046
rect 7786 2810 8022 3046
rect 9286 28310 9522 28546
rect 9286 25536 9316 25546
rect 9316 25536 9332 25546
rect 9332 25536 9396 25546
rect 9396 25536 9412 25546
rect 9412 25536 9476 25546
rect 9476 25536 9492 25546
rect 9492 25536 9522 25546
rect 9286 25310 9522 25536
rect 9286 22336 9522 22546
rect 9286 22310 9316 22336
rect 9316 22310 9332 22336
rect 9332 22310 9396 22336
rect 9396 22310 9412 22336
rect 9412 22310 9476 22336
rect 9476 22310 9492 22336
rect 9492 22310 9522 22336
rect 9286 19310 9522 19546
rect 9286 16310 9522 16546
rect 9286 13310 9522 13546
rect 9286 10368 9522 10546
rect 9286 10310 9316 10368
rect 9316 10310 9332 10368
rect 9332 10310 9396 10368
rect 9396 10310 9412 10368
rect 9412 10310 9476 10368
rect 9476 10310 9492 10368
rect 9492 10310 9522 10368
rect 9286 7310 9522 7546
rect 9286 4310 9522 4546
rect 10786 26810 11022 27046
rect 10786 23968 11022 24046
rect 10786 23904 10816 23968
rect 10816 23904 10832 23968
rect 10832 23904 10896 23968
rect 10896 23904 10912 23968
rect 10912 23904 10976 23968
rect 10976 23904 10992 23968
rect 10992 23904 11022 23968
rect 10786 23810 11022 23904
rect 10786 20810 11022 21046
rect 10786 17810 11022 18046
rect 10786 14810 11022 15046
rect 10786 12000 11022 12046
rect 10786 11936 10816 12000
rect 10816 11936 10832 12000
rect 10832 11936 10896 12000
rect 10896 11936 10912 12000
rect 10912 11936 10976 12000
rect 10976 11936 10992 12000
rect 10992 11936 11022 12000
rect 10786 11810 11022 11936
rect 10786 8810 11022 9046
rect 10786 5810 11022 6046
rect 10786 2810 11022 3046
rect 12286 28310 12522 28546
rect 12286 25536 12316 25546
rect 12316 25536 12332 25546
rect 12332 25536 12396 25546
rect 12396 25536 12412 25546
rect 12412 25536 12476 25546
rect 12476 25536 12492 25546
rect 12492 25536 12522 25546
rect 12286 25310 12522 25536
rect 12286 22336 12522 22546
rect 12286 22310 12316 22336
rect 12316 22310 12332 22336
rect 12332 22310 12396 22336
rect 12396 22310 12412 22336
rect 12412 22310 12476 22336
rect 12476 22310 12492 22336
rect 12492 22310 12522 22336
rect 12286 19310 12522 19546
rect 12286 16310 12522 16546
rect 12286 13310 12522 13546
rect 12286 10368 12522 10546
rect 12286 10310 12316 10368
rect 12316 10310 12332 10368
rect 12332 10310 12396 10368
rect 12396 10310 12412 10368
rect 12412 10310 12476 10368
rect 12476 10310 12492 10368
rect 12492 10310 12522 10368
rect 12286 7310 12522 7546
rect 12286 4310 12522 4546
rect 13786 26810 14022 27046
rect 13786 23968 14022 24046
rect 13786 23904 13816 23968
rect 13816 23904 13832 23968
rect 13832 23904 13896 23968
rect 13896 23904 13912 23968
rect 13912 23904 13976 23968
rect 13976 23904 13992 23968
rect 13992 23904 14022 23968
rect 13786 23810 14022 23904
rect 13786 20810 14022 21046
rect 13786 17810 14022 18046
rect 13786 14810 14022 15046
rect 13786 12000 14022 12046
rect 13786 11936 13816 12000
rect 13816 11936 13832 12000
rect 13832 11936 13896 12000
rect 13896 11936 13912 12000
rect 13912 11936 13976 12000
rect 13976 11936 13992 12000
rect 13992 11936 14022 12000
rect 13786 11810 14022 11936
rect 13786 8810 14022 9046
rect 13786 5810 14022 6046
rect 13786 2810 14022 3046
rect 15286 28310 15522 28546
rect 15286 25536 15316 25546
rect 15316 25536 15332 25546
rect 15332 25536 15396 25546
rect 15396 25536 15412 25546
rect 15412 25536 15476 25546
rect 15476 25536 15492 25546
rect 15492 25536 15522 25546
rect 15286 25310 15522 25536
rect 15286 22336 15522 22546
rect 15286 22310 15316 22336
rect 15316 22310 15332 22336
rect 15332 22310 15396 22336
rect 15396 22310 15412 22336
rect 15412 22310 15476 22336
rect 15476 22310 15492 22336
rect 15492 22310 15522 22336
rect 15286 19310 15522 19546
rect 15286 16310 15522 16546
rect 15286 13310 15522 13546
rect 15286 10368 15522 10546
rect 15286 10310 15316 10368
rect 15316 10310 15332 10368
rect 15332 10310 15396 10368
rect 15396 10310 15412 10368
rect 15412 10310 15476 10368
rect 15476 10310 15492 10368
rect 15492 10310 15522 10368
rect 15286 7310 15522 7546
rect 15286 4310 15522 4546
rect 16786 26810 17022 27046
rect 16786 23968 17022 24046
rect 16786 23904 16816 23968
rect 16816 23904 16832 23968
rect 16832 23904 16896 23968
rect 16896 23904 16912 23968
rect 16912 23904 16976 23968
rect 16976 23904 16992 23968
rect 16992 23904 17022 23968
rect 16786 23810 17022 23904
rect 16786 20810 17022 21046
rect 16786 17810 17022 18046
rect 16786 14810 17022 15046
rect 16786 12000 17022 12046
rect 16786 11936 16816 12000
rect 16816 11936 16832 12000
rect 16832 11936 16896 12000
rect 16896 11936 16912 12000
rect 16912 11936 16976 12000
rect 16976 11936 16992 12000
rect 16992 11936 17022 12000
rect 16786 11810 17022 11936
rect 16786 8810 17022 9046
rect 16786 5810 17022 6046
rect 16786 2810 17022 3046
rect 18286 28310 18522 28546
rect 18286 25536 18316 25546
rect 18316 25536 18332 25546
rect 18332 25536 18396 25546
rect 18396 25536 18412 25546
rect 18412 25536 18476 25546
rect 18476 25536 18492 25546
rect 18492 25536 18522 25546
rect 18286 25310 18522 25536
rect 18286 22336 18522 22546
rect 18286 22310 18316 22336
rect 18316 22310 18332 22336
rect 18332 22310 18396 22336
rect 18396 22310 18412 22336
rect 18412 22310 18476 22336
rect 18476 22310 18492 22336
rect 18492 22310 18522 22336
rect 18286 19310 18522 19546
rect 18286 16310 18522 16546
rect 18286 13310 18522 13546
rect 18286 10368 18522 10546
rect 18286 10310 18316 10368
rect 18316 10310 18332 10368
rect 18332 10310 18396 10368
rect 18396 10310 18412 10368
rect 18412 10310 18476 10368
rect 18476 10310 18492 10368
rect 18492 10310 18522 10368
rect 18286 7310 18522 7546
rect 18286 4310 18522 4546
rect 19786 26810 20022 27046
rect 19786 23968 20022 24046
rect 19786 23904 19816 23968
rect 19816 23904 19832 23968
rect 19832 23904 19896 23968
rect 19896 23904 19912 23968
rect 19912 23904 19976 23968
rect 19976 23904 19992 23968
rect 19992 23904 20022 23968
rect 19786 23810 20022 23904
rect 19786 20810 20022 21046
rect 19786 17810 20022 18046
rect 19786 14810 20022 15046
rect 19786 12000 20022 12046
rect 19786 11936 19816 12000
rect 19816 11936 19832 12000
rect 19832 11936 19896 12000
rect 19896 11936 19912 12000
rect 19912 11936 19976 12000
rect 19976 11936 19992 12000
rect 19992 11936 20022 12000
rect 19786 11810 20022 11936
rect 19786 8810 20022 9046
rect 19786 5810 20022 6046
rect 19786 2810 20022 3046
rect 21286 28310 21522 28546
rect 21286 25536 21316 25546
rect 21316 25536 21332 25546
rect 21332 25536 21396 25546
rect 21396 25536 21412 25546
rect 21412 25536 21476 25546
rect 21476 25536 21492 25546
rect 21492 25536 21522 25546
rect 21286 25310 21522 25536
rect 21286 22336 21522 22546
rect 21286 22310 21316 22336
rect 21316 22310 21332 22336
rect 21332 22310 21396 22336
rect 21396 22310 21412 22336
rect 21412 22310 21476 22336
rect 21476 22310 21492 22336
rect 21492 22310 21522 22336
rect 21286 19310 21522 19546
rect 21286 16310 21522 16546
rect 21286 13310 21522 13546
rect 21286 10368 21522 10546
rect 21286 10310 21316 10368
rect 21316 10310 21332 10368
rect 21332 10310 21396 10368
rect 21396 10310 21412 10368
rect 21412 10310 21476 10368
rect 21476 10310 21492 10368
rect 21492 10310 21522 10368
rect 21286 7310 21522 7546
rect 21286 4310 21522 4546
rect 22786 26810 23022 27046
rect 22786 23968 23022 24046
rect 22786 23904 22816 23968
rect 22816 23904 22832 23968
rect 22832 23904 22896 23968
rect 22896 23904 22912 23968
rect 22912 23904 22976 23968
rect 22976 23904 22992 23968
rect 22992 23904 23022 23968
rect 22786 23810 23022 23904
rect 22786 20810 23022 21046
rect 22786 17810 23022 18046
rect 22786 14810 23022 15046
rect 22786 12000 23022 12046
rect 22786 11936 22816 12000
rect 22816 11936 22832 12000
rect 22832 11936 22896 12000
rect 22896 11936 22912 12000
rect 22912 11936 22976 12000
rect 22976 11936 22992 12000
rect 22992 11936 23022 12000
rect 22786 11810 23022 11936
rect 22786 8810 23022 9046
rect 22786 5810 23022 6046
rect 22786 2810 23022 3046
rect 24286 28310 24522 28546
rect 24286 25536 24316 25546
rect 24316 25536 24332 25546
rect 24332 25536 24396 25546
rect 24396 25536 24412 25546
rect 24412 25536 24476 25546
rect 24476 25536 24492 25546
rect 24492 25536 24522 25546
rect 24286 25310 24522 25536
rect 24286 22336 24522 22546
rect 24286 22310 24316 22336
rect 24316 22310 24332 22336
rect 24332 22310 24396 22336
rect 24396 22310 24412 22336
rect 24412 22310 24476 22336
rect 24476 22310 24492 22336
rect 24492 22310 24522 22336
rect 24286 19310 24522 19546
rect 24286 16310 24522 16546
rect 24286 13310 24522 13546
rect 24286 10368 24522 10546
rect 24286 10310 24316 10368
rect 24316 10310 24332 10368
rect 24332 10310 24396 10368
rect 24396 10310 24412 10368
rect 24412 10310 24476 10368
rect 24476 10310 24492 10368
rect 24492 10310 24522 10368
rect 24286 7310 24522 7546
rect 24286 4310 24522 4546
rect 25786 26810 26022 27046
rect 25786 23968 26022 24046
rect 25786 23904 25816 23968
rect 25816 23904 25832 23968
rect 25832 23904 25896 23968
rect 25896 23904 25912 23968
rect 25912 23904 25976 23968
rect 25976 23904 25992 23968
rect 25992 23904 26022 23968
rect 25786 23810 26022 23904
rect 25786 20810 26022 21046
rect 25786 17810 26022 18046
rect 25786 14810 26022 15046
rect 25786 12000 26022 12046
rect 25786 11936 25816 12000
rect 25816 11936 25832 12000
rect 25832 11936 25896 12000
rect 25896 11936 25912 12000
rect 25912 11936 25976 12000
rect 25976 11936 25992 12000
rect 25992 11936 26022 12000
rect 25786 11810 26022 11936
rect 25786 8810 26022 9046
rect 25786 5810 26022 6046
rect 25786 2810 26022 3046
rect 27286 28310 27522 28546
rect 27286 25536 27316 25546
rect 27316 25536 27332 25546
rect 27332 25536 27396 25546
rect 27396 25536 27412 25546
rect 27412 25536 27476 25546
rect 27476 25536 27492 25546
rect 27492 25536 27522 25546
rect 27286 25310 27522 25536
rect 27286 22336 27522 22546
rect 27286 22310 27316 22336
rect 27316 22310 27332 22336
rect 27332 22310 27396 22336
rect 27396 22310 27412 22336
rect 27412 22310 27476 22336
rect 27476 22310 27492 22336
rect 27492 22310 27522 22336
rect 27286 19310 27522 19546
rect 27286 16310 27522 16546
rect 27286 13310 27522 13546
rect 27286 10368 27522 10546
rect 27286 10310 27316 10368
rect 27316 10310 27332 10368
rect 27332 10310 27396 10368
rect 27396 10310 27412 10368
rect 27412 10310 27476 10368
rect 27476 10310 27492 10368
rect 27492 10310 27522 10368
rect 27286 7310 27522 7546
rect 27286 4310 27522 4546
<< metal5 >>
rect 1104 28546 28336 28588
rect 1104 28310 3286 28546
rect 3522 28310 6286 28546
rect 6522 28310 9286 28546
rect 9522 28310 12286 28546
rect 12522 28310 15286 28546
rect 15522 28310 18286 28546
rect 18522 28310 21286 28546
rect 21522 28310 24286 28546
rect 24522 28310 27286 28546
rect 27522 28310 28336 28546
rect 1104 28268 28336 28310
rect 1104 27046 28336 27088
rect 1104 26810 1786 27046
rect 2022 26810 4786 27046
rect 5022 26810 7786 27046
rect 8022 26810 10786 27046
rect 11022 26810 13786 27046
rect 14022 26810 16786 27046
rect 17022 26810 19786 27046
rect 20022 26810 22786 27046
rect 23022 26810 25786 27046
rect 26022 26810 28336 27046
rect 1104 26768 28336 26810
rect 1104 25546 28336 25588
rect 1104 25310 3286 25546
rect 3522 25310 6286 25546
rect 6522 25310 9286 25546
rect 9522 25310 12286 25546
rect 12522 25310 15286 25546
rect 15522 25310 18286 25546
rect 18522 25310 21286 25546
rect 21522 25310 24286 25546
rect 24522 25310 27286 25546
rect 27522 25310 28336 25546
rect 1104 25268 28336 25310
rect 1104 24046 28336 24088
rect 1104 23810 1786 24046
rect 2022 23810 4786 24046
rect 5022 23810 7786 24046
rect 8022 23810 10786 24046
rect 11022 23810 13786 24046
rect 14022 23810 16786 24046
rect 17022 23810 19786 24046
rect 20022 23810 22786 24046
rect 23022 23810 25786 24046
rect 26022 23810 28336 24046
rect 1104 23768 28336 23810
rect 1104 22546 28336 22588
rect 1104 22310 3286 22546
rect 3522 22310 6286 22546
rect 6522 22310 9286 22546
rect 9522 22310 12286 22546
rect 12522 22310 15286 22546
rect 15522 22310 18286 22546
rect 18522 22310 21286 22546
rect 21522 22310 24286 22546
rect 24522 22310 27286 22546
rect 27522 22310 28336 22546
rect 1104 22268 28336 22310
rect 1104 21046 28336 21088
rect 1104 20810 1786 21046
rect 2022 20810 4786 21046
rect 5022 20810 7786 21046
rect 8022 20810 10786 21046
rect 11022 20810 13786 21046
rect 14022 20810 16786 21046
rect 17022 20810 19786 21046
rect 20022 20810 22786 21046
rect 23022 20810 25786 21046
rect 26022 20810 28336 21046
rect 1104 20768 28336 20810
rect 1104 19546 28336 19588
rect 1104 19310 3286 19546
rect 3522 19310 6286 19546
rect 6522 19310 9286 19546
rect 9522 19310 12286 19546
rect 12522 19310 15286 19546
rect 15522 19310 18286 19546
rect 18522 19310 21286 19546
rect 21522 19310 24286 19546
rect 24522 19310 27286 19546
rect 27522 19310 28336 19546
rect 1104 19268 28336 19310
rect 1104 18046 28336 18088
rect 1104 17810 1786 18046
rect 2022 17810 4786 18046
rect 5022 17810 7786 18046
rect 8022 17810 10786 18046
rect 11022 17810 13786 18046
rect 14022 17810 16786 18046
rect 17022 17810 19786 18046
rect 20022 17810 22786 18046
rect 23022 17810 25786 18046
rect 26022 17810 28336 18046
rect 1104 17768 28336 17810
rect 1104 16546 28336 16588
rect 1104 16310 3286 16546
rect 3522 16310 6286 16546
rect 6522 16310 9286 16546
rect 9522 16310 12286 16546
rect 12522 16310 15286 16546
rect 15522 16310 18286 16546
rect 18522 16310 21286 16546
rect 21522 16310 24286 16546
rect 24522 16310 27286 16546
rect 27522 16310 28336 16546
rect 1104 16268 28336 16310
rect 1104 15046 28336 15088
rect 1104 14810 1786 15046
rect 2022 14810 4786 15046
rect 5022 14810 7786 15046
rect 8022 14810 10786 15046
rect 11022 14810 13786 15046
rect 14022 14810 16786 15046
rect 17022 14810 19786 15046
rect 20022 14810 22786 15046
rect 23022 14810 25786 15046
rect 26022 14810 28336 15046
rect 1104 14768 28336 14810
rect 1104 13546 28336 13588
rect 1104 13310 3286 13546
rect 3522 13310 6286 13546
rect 6522 13310 9286 13546
rect 9522 13310 12286 13546
rect 12522 13310 15286 13546
rect 15522 13310 18286 13546
rect 18522 13310 21286 13546
rect 21522 13310 24286 13546
rect 24522 13310 27286 13546
rect 27522 13310 28336 13546
rect 1104 13268 28336 13310
rect 1104 12046 28336 12088
rect 1104 11810 1786 12046
rect 2022 11810 4786 12046
rect 5022 11810 7786 12046
rect 8022 11810 10786 12046
rect 11022 11810 13786 12046
rect 14022 11810 16786 12046
rect 17022 11810 19786 12046
rect 20022 11810 22786 12046
rect 23022 11810 25786 12046
rect 26022 11810 28336 12046
rect 1104 11768 28336 11810
rect 1104 10546 28336 10588
rect 1104 10310 3286 10546
rect 3522 10310 6286 10546
rect 6522 10310 9286 10546
rect 9522 10310 12286 10546
rect 12522 10310 15286 10546
rect 15522 10310 18286 10546
rect 18522 10310 21286 10546
rect 21522 10310 24286 10546
rect 24522 10310 27286 10546
rect 27522 10310 28336 10546
rect 1104 10268 28336 10310
rect 1104 9046 28336 9088
rect 1104 8810 1786 9046
rect 2022 8810 4786 9046
rect 5022 8810 7786 9046
rect 8022 8810 10786 9046
rect 11022 8810 13786 9046
rect 14022 8810 16786 9046
rect 17022 8810 19786 9046
rect 20022 8810 22786 9046
rect 23022 8810 25786 9046
rect 26022 8810 28336 9046
rect 1104 8768 28336 8810
rect 1104 7546 28336 7588
rect 1104 7310 3286 7546
rect 3522 7310 6286 7546
rect 6522 7310 9286 7546
rect 9522 7310 12286 7546
rect 12522 7310 15286 7546
rect 15522 7310 18286 7546
rect 18522 7310 21286 7546
rect 21522 7310 24286 7546
rect 24522 7310 27286 7546
rect 27522 7310 28336 7546
rect 1104 7268 28336 7310
rect 1104 6046 28336 6088
rect 1104 5810 1786 6046
rect 2022 5810 4786 6046
rect 5022 5810 7786 6046
rect 8022 5810 10786 6046
rect 11022 5810 13786 6046
rect 14022 5810 16786 6046
rect 17022 5810 19786 6046
rect 20022 5810 22786 6046
rect 23022 5810 25786 6046
rect 26022 5810 28336 6046
rect 1104 5768 28336 5810
rect 1104 4546 28336 4588
rect 1104 4310 3286 4546
rect 3522 4310 6286 4546
rect 6522 4310 9286 4546
rect 9522 4310 12286 4546
rect 12522 4310 15286 4546
rect 15522 4310 18286 4546
rect 18522 4310 21286 4546
rect 21522 4310 24286 4546
rect 24522 4310 27286 4546
rect 27522 4310 28336 4546
rect 1104 4268 28336 4310
rect 1104 3046 28336 3088
rect 1104 2810 1786 3046
rect 2022 2810 4786 3046
rect 5022 2810 7786 3046
rect 8022 2810 10786 3046
rect 11022 2810 13786 3046
rect 14022 2810 16786 3046
rect 17022 2810 19786 3046
rect 20022 2810 22786 3046
rect 23022 2810 25786 3046
rect 26022 2810 28336 3046
rect 1104 2768 28336 2810
use sky130_fd_sc_hd__decap_12  FILLER_2_15 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1597341371
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1597341371
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1597341371
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1597341371
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1597341371
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1597341371
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1597341371
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1597341371
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1597341371
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1597341371
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1597341371
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1597341371
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1597341371
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1597341371
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1597341371
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_62 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_56 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1597341371
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1597341371
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1597341371
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A1 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1597341371
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1597341371
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1597341371
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1597341371
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1597341371
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A1
timestamp 1597341371
transform 1 0 6900 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1597341371
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1597341371
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1597341371
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1597341371
transform 1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1597341371
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__B1_N
timestamp 1597341371
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _148_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74
timestamp 1597341371
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1597341371
transform 1 0 7820 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A2
timestamp 1597341371
transform 1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _206_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7636 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1597341371
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__D
timestamp 1597341371
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1597341371
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1597341371
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__RESET_B
timestamp 1597341371
transform 1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__RESET_B
timestamp 1597341371
transform 1 0 8556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1597341371
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_84
timestamp 1597341371
transform 1 0 8832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1597341371
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__D
timestamp 1597341371
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__CLK
timestamp 1597341371
transform 1 0 9016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1597341371
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1597341371
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1597341371
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1597341371
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1597341371
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__CLK
timestamp 1597341371
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1597341371
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1597341371
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1597341371
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1597341371
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp 1597341371
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1597341371
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1597341371
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__B1
timestamp 1597341371
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _290_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 9476 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1597341371
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1597341371
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A2
timestamp 1597341371
transform 1 0 10396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__B
timestamp 1597341371
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _201_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 11132 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_2_113
timestamp 1597341371
transform 1 0 11500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_114
timestamp 1597341371
transform 1 0 11592 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_116
timestamp 1597341371
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A1
timestamp 1597341371
transform 1 0 11776 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1597341371
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1597341371
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__B1
timestamp 1597341371
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A2
timestamp 1597341371
transform 1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__RESET_B
timestamp 1597341371
transform 1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_122
timestamp 1597341371
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1597341371
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1597341371
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1597341371
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1597341371
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _204_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _202_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 12512 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1597341371
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134
timestamp 1597341371
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_130
timestamp 1597341371
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1597341371
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__D
timestamp 1597341371
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__CLK
timestamp 1597341371
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1597341371
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1597341371
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1597341371
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1597341371
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_147
timestamp 1597341371
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1597341371
transform 1 0 14628 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__C
timestamp 1597341371
transform 1 0 13892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__C
timestamp 1597341371
transform 1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _203_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 13800 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _289_
timestamp 1597341371
transform 1 0 12880 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1597341371
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1597341371
transform 1 0 14996 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1597341371
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1597341371
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__D
timestamp 1597341371
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1597341371
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1597341371
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1597341371
transform 1 0 15640 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_161
timestamp 1597341371
transform 1 0 15916 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157
timestamp 1597341371
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1597341371
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__CLK
timestamp 1597341371
transform 1 0 15732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _200_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15640 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_165
timestamp 1597341371
transform 1 0 16284 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_171
timestamp 1597341371
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_167
timestamp 1597341371
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__B
timestamp 1597341371
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1597341371
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _140_
timestamp 1597341371
transform 1 0 16376 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_4  _278_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15732 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1597341371
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1597341371
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 1597341371
transform 1 0 17388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__SET_B
timestamp 1597341371
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1597341371
transform 1 0 17940 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1597341371
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_179
timestamp 1597341371
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1597341371
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1597341371
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1597341371
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1597341371
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__C
timestamp 1597341371
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1597341371
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1597341371
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_187
timestamp 1597341371
transform 1 0 18308 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1597341371
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1597341371
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1597341371
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1597341371
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _146_
timestamp 1597341371
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1597341371
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1597341371
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1597341371
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1597341371
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_198
timestamp 1597341371
transform 1 0 19320 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1597341371
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__D
timestamp 1597341371
transform 1 0 19136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1597341371
transform 1 0 19136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_198
timestamp 1597341371
transform 1 0 19320 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_207
timestamp 1597341371
transform 1 0 20148 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1597341371
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_210
timestamp 1597341371
transform 1 0 20424 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__B
timestamp 1597341371
transform 1 0 19964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1597341371
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1597341371
transform 1 0 19596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1597341371
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1597341371
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1597341371
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1597341371
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1597341371
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_213
timestamp 1597341371
transform 1 0 20700 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_201
timestamp 1597341371
transform 1 0 19596 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1597341371
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1597341371
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1597341371
transform 1 0 22908 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1597341371
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1597341371
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1597341371
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1597341371
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1597341371
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1597341371
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1597341371
transform 1 0 21804 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1597341371
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1597341371
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1597341371
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1597341371
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1597341371
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1597341371
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1597341371
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1597341371
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1597341371
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1597341371
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_292
timestamp 1597341371
transform 1 0 27968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_288
timestamp 1597341371
transform 1 0 27600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_292
timestamp 1597341371
transform 1 0 27968 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1597341371
transform -1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1597341371
transform -1 0 28336 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1597341371
transform -1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1597341371
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1597341371
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1597341371
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1597341371
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1597341371
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1597341371
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1597341371
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1597341371
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1597341371
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1597341371
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1597341371
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1597341371
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1597341371
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1597341371
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1597341371
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1597341371
transform 1 0 6256 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1597341371
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1597341371
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_60
timestamp 1597341371
transform 1 0 6624 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1597341371
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1597341371
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1597341371
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1597341371
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1597341371
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1597341371
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1597341371
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B2
timestamp 1597341371
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__B1
timestamp 1597341371
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A2
timestamp 1597341371
transform 1 0 7544 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B1
timestamp 1597341371
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1597341371
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1597341371
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A2
timestamp 1597341371
transform 1 0 7820 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__B
timestamp 1597341371
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1597341371
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1597341371
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp 1597341371
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__B1
timestamp 1597341371
transform 1 0 9016 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _205_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_4_98
timestamp 1597341371
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1597341371
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1597341371
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__C
timestamp 1597341371
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1597341371
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _291_
timestamp 1597341371
transform 1 0 8280 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_3_109
timestamp 1597341371
transform 1 0 11132 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_105
timestamp 1597341371
transform 1 0 10764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1597341371
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__B
timestamp 1597341371
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A1
timestamp 1597341371
transform 1 0 10580 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1597341371
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_116
timestamp 1597341371
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1597341371
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1597341371
transform 1 0 11592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__B
timestamp 1597341371
transform 1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1597341371
transform 1 0 11960 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1597341371
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1597341371
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__C
timestamp 1597341371
transform 1 0 11960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1597341371
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _167_
timestamp 1597341371
transform 1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _169_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 10304 0 1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_4_131
timestamp 1597341371
transform 1 0 13156 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1597341371
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _166_
timestamp 1597341371
transform 1 0 12696 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_140
timestamp 1597341371
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_136
timestamp 1597341371
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1597341371
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1597341371
transform 1 0 13524 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1597341371
transform 1 0 13892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__B1
timestamp 1597341371
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _195_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 14260 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1597341371
transform 1 0 14168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1597341371
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1597341371
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1597341371
transform 1 0 14628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1597341371
transform 1 0 15640 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1597341371
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_161
timestamp 1597341371
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1597341371
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_152
timestamp 1597341371
transform 1 0 15088 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__D
timestamp 1597341371
transform 1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__CLK
timestamp 1597341371
transform 1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1597341371
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1597341371
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _173_
timestamp 1597341371
transform 1 0 16100 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _279_
timestamp 1597341371
transform 1 0 15732 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1597341371
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1597341371
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_176
timestamp 1597341371
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1597341371
transform 1 0 17480 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__RESET_B
timestamp 1597341371
transform 1 0 17112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1597341371
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1597341371
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1597341371
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1597341371
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__D
timestamp 1597341371
transform 1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _199_
timestamp 1597341371
transform 1 0 18216 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp 1597341371
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1597341371
transform 1 0 19228 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1597341371
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__RESET_B
timestamp 1597341371
transform 1 0 19228 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__CLK
timestamp 1597341371
transform 1 0 19044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_199
timestamp 1597341371
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1597341371
transform 1 0 19596 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1597341371
transform 1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1597341371
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1597341371
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1597341371
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1597341371
transform 1 0 20056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_208
timestamp 1597341371
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1597341371
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1597341371
transform 1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1597341371
transform 1 0 20424 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_219
timestamp 1597341371
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1597341371
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1597341371
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A1
timestamp 1597341371
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B2
timestamp 1597341371
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1597341371
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_223
timestamp 1597341371
transform 1 0 21620 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_212
timestamp 1597341371
transform 1 0 20608 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_247
timestamp 1597341371
transform 1 0 23828 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_235
timestamp 1597341371
transform 1 0 22724 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1597341371
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_236 home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 22816 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_224
timestamp 1597341371
transform 1 0 21712 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1597341371
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1597341371
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1597341371
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1597341371
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1597341371
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_292
timestamp 1597341371
transform 1 0 27968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1597341371
transform 1 0 27600 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1597341371
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1597341371
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1597341371
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1597341371
transform -1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1597341371
transform -1 0 28336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1597341371
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1597341371
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1597341371
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1597341371
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1597341371
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1597341371
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1597341371
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_44
timestamp 1597341371
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1597341371
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1597341371
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1597341371
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1597341371
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__B
timestamp 1597341371
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1597341371
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_52
timestamp 1597341371
transform 1 0 5888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__A
timestamp 1597341371
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1597341371
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1597341371
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1597341371
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1597341371
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B2
timestamp 1597341371
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__RESET_B
timestamp 1597341371
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1597341371
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1597341371
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 1597341371
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1597341371
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1597341371
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A1
timestamp 1597341371
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__D
timestamp 1597341371
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__293__CLK
timestamp 1597341371
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _293_
timestamp 1597341371
transform 1 0 6716 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1597341371
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1597341371
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A3
timestamp 1597341371
transform 1 0 9016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A2
timestamp 1597341371
transform 1 0 8096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1597341371
transform 1 0 10028 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1597341371
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1597341371
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1597341371
transform 1 0 9752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1597341371
transform 1 0 10120 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A
timestamp 1597341371
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1597341371
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _275_
timestamp 1597341371
transform 1 0 8648 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_108
timestamp 1597341371
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_104
timestamp 1597341371
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1597341371
transform 1 0 10396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1597341371
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__B
timestamp 1597341371
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1597341371
transform 1 0 10856 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _165_
timestamp 1597341371
transform 1 0 10488 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_119
timestamp 1597341371
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1597341371
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1597341371
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_111
timestamp 1597341371
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1597341371
transform 1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__D
timestamp 1597341371
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _196_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 11224 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1597341371
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A2
timestamp 1597341371
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1597341371
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_134
timestamp 1597341371
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1597341371
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_134
timestamp 1597341371
transform 1 0 13432 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _178_
timestamp 1597341371
transform 1 0 12604 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _168_
timestamp 1597341371
transform 1 0 12788 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_138
timestamp 1597341371
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1597341371
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1597341371
transform 1 0 13800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__C1
timestamp 1597341371
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B1
timestamp 1597341371
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1597341371
transform 1 0 14168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1597341371
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1597341371
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1597341371
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__B
timestamp 1597341371
transform 1 0 14628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _179_
timestamp 1597341371
transform 1 0 14536 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1597341371
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_159
timestamp 1597341371
transform 1 0 15732 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1597341371
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A2
timestamp 1597341371
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1597341371
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1597341371
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1597341371
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B
timestamp 1597341371
transform 1 0 16928 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__B1
timestamp 1597341371
transform 1 0 16928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _180_
timestamp 1597341371
transform 1 0 16100 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _270_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15456 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_6_178
timestamp 1597341371
transform 1 0 17480 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1597341371
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1597341371
transform 1 0 17480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1597341371
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A2
timestamp 1597341371
transform 1 0 17296 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A1
timestamp 1597341371
transform 1 0 17296 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1597341371
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1597341371
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _221_
timestamp 1597341371
transform 1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_184
timestamp 1597341371
transform 1 0 18032 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1597341371
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1597341371
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1597341371
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_188
timestamp 1597341371
transform 1 0 18400 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A2
timestamp 1597341371
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _216_
timestamp 1597341371
transform 1 0 18768 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  _281_
timestamp 1597341371
transform 1 0 18676 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_6_208
timestamp 1597341371
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp 1597341371
transform 1 0 19780 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_199
timestamp 1597341371
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 1597341371
transform 1 0 19596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__D
timestamp 1597341371
transform 1 0 20056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__CLK
timestamp 1597341371
transform 1 0 20424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1597341371
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1597341371
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1597341371
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1597341371
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_214
timestamp 1597341371
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A2
timestamp 1597341371
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__RESET_B
timestamp 1597341371
transform 1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1597341371
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _223_
timestamp 1597341371
transform 1 0 21068 0 1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_6_243
timestamp 1597341371
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_231
timestamp 1597341371
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1597341371
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_238
timestamp 1597341371
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_226
timestamp 1597341371
transform 1 0 21896 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__B1
timestamp 1597341371
transform 1 0 21712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1597341371
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_267
timestamp 1597341371
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_255
timestamp 1597341371
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1597341371
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1597341371
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_292
timestamp 1597341371
transform 1 0 27968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1597341371
transform 1 0 27600 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1597341371
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1597341371
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1597341371
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1597341371
transform -1 0 28336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1597341371
transform -1 0 28336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1597341371
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1597341371
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1597341371
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1597341371
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1597341371
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1597341371
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1597341371
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1597341371
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1597341371
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_45
timestamp 1597341371
transform 1 0 5244 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_39
timestamp 1597341371
transform 1 0 4692 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1597341371
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1597341371
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _272_
timestamp 1597341371
transform 1 0 5336 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_59
timestamp 1597341371
transform 1 0 6532 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1597341371
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1597341371
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1597341371
transform 1 0 5980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1597341371
transform 1 0 6256 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1597341371
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1597341371
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1597341371
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_67
timestamp 1597341371
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A
timestamp 1597341371
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__B
timestamp 1597341371
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _273_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7268 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _276_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 7452 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_8_84
timestamp 1597341371
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1597341371
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp 1597341371
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1597341371
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__B
timestamp 1597341371
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1597341371
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1597341371
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1597341371
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1597341371
transform 1 0 9016 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B
timestamp 1597341371
transform 1 0 9200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A
timestamp 1597341371
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1597341371
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _274_
timestamp 1597341371
transform 1 0 9752 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _171_
timestamp 1597341371
transform 1 0 9844 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1597341371
transform 1 0 11040 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1597341371
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1597341371
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_105
timestamp 1597341371
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1597341371
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1597341371
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__RESET_B
timestamp 1597341371
transform 1 0 10580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__D
timestamp 1597341371
transform 1 0 10948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp 1597341371
transform 1 0 11316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1597341371
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1597341371
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1597341371
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__CLK
timestamp 1597341371
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1597341371
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _292_
timestamp 1597341371
transform 1 0 11408 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_8_135
timestamp 1597341371
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_139
timestamp 1597341371
transform 1 0 13892 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1597341371
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_137
timestamp 1597341371
transform 1 0 13708 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__B
timestamp 1597341371
transform 1 0 13984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A2_N
timestamp 1597341371
transform 1 0 14168 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1597341371
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1597341371
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1597341371
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A1_N
timestamp 1597341371
transform 1 0 14536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _269_
timestamp 1597341371
transform 1 0 14352 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _197_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1597341371
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1597341371
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_159
timestamp 1597341371
transform 1 0 15732 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1597341371
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1597341371
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1597341371
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1597341371
transform 1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1597341371
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _213_
timestamp 1597341371
transform 1 0 15456 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_172
timestamp 1597341371
transform 1 0 16928 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_167
timestamp 1597341371
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1597341371
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B2
timestamp 1597341371
transform 1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1597341371
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _214_
timestamp 1597341371
transform 1 0 16100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_183
timestamp 1597341371
transform 1 0 17940 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp 1597341371
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1597341371
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1597341371
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1597341371
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1597341371
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1597341371
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _160_
timestamp 1597341371
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_195
timestamp 1597341371
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_191
timestamp 1597341371
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_187
timestamp 1597341371
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1597341371
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B
timestamp 1597341371
transform 1 0 18492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1597341371
transform 1 0 18860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__B2
timestamp 1597341371
transform 1 0 18308 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _207_
timestamp 1597341371
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _215_
timestamp 1597341371
transform 1 0 18676 0 -1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1597341371
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1597341371
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1597341371
transform 1 0 20332 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_205
timestamp 1597341371
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1597341371
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A1
timestamp 1597341371
transform 1 0 20148 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_219
timestamp 1597341371
transform 1 0 21252 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1597341371
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A2
timestamp 1597341371
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1597341371
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1597341371
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _282_
timestamp 1597341371
transform 1 0 20700 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_8_244
timestamp 1597341371
transform 1 0 23552 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_232
timestamp 1597341371
transform 1 0 22448 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_228
timestamp 1597341371
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_224
timestamp 1597341371
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1597341371
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_236
timestamp 1597341371
transform 1 0 22816 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1597341371
transform 1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1597341371
transform 1 0 21896 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1597341371
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_268
timestamp 1597341371
transform 1 0 25760 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_256
timestamp 1597341371
transform 1 0 24656 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1597341371
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1597341371
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_292
timestamp 1597341371
transform 1 0 27968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1597341371
transform 1 0 27600 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1597341371
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1597341371
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1597341371
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1597341371
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1597341371
transform -1 0 28336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1597341371
transform -1 0 28336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1597341371
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1597341371
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1597341371
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1597341371
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1597341371
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1597341371
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1597341371
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1597341371
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1597341371
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1597341371
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1597341371
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1597341371
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1597341371
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_56
timestamp 1597341371
transform 1 0 6256 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1597341371
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1597341371
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1597341371
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A1
timestamp 1597341371
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__B
timestamp 1597341371
transform 1 0 6716 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1597341371
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_63
timestamp 1597341371
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1597341371
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A2
timestamp 1597341371
transform 1 0 6992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1597341371
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1597341371
transform 1 0 7636 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1597341371
transform 1 0 7268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1597341371
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A1
timestamp 1597341371
transform 1 0 7360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1597341371
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__B1
timestamp 1597341371
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _271_
timestamp 1597341371
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1597341371
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1597341371
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A2
timestamp 1597341371
transform 1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _177_
timestamp 1597341371
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1597341371
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1597341371
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1597341371
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B1
timestamp 1597341371
transform 1 0 9016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__B
timestamp 1597341371
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1597341371
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_99
timestamp 1597341371
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1597341371
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B
timestamp 1597341371
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _208_
timestamp 1597341371
transform 1 0 9844 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1597341371
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 1597341371
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1597341371
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1597341371
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1597341371
transform 1 0 11040 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 1597341371
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1597341371
transform 1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_112
timestamp 1597341371
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1597341371
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1597341371
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1597341371
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_116
timestamp 1597341371
transform 1 0 11776 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1597341371
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__C
timestamp 1597341371
transform 1 0 11592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1597341371
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1597341371
transform 1 0 11960 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1597341371
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1597341371
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1597341371
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__CLK
timestamp 1597341371
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1597341371
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__RESET_B
timestamp 1597341371
transform 1 0 12512 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1597341371
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_130
timestamp 1597341371
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1597341371
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1597341371
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1597341371
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__D
timestamp 1597341371
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1597341371
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _139_
timestamp 1597341371
transform 1 0 12604 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1597341371
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1597341371
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1597341371
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_138
timestamp 1597341371
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 1597341371
transform 1 0 14168 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A
timestamp 1597341371
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__B1
timestamp 1597341371
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _268_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 14536 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1597341371
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1597341371
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1597341371
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1597341371
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 1597341371
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_161
timestamp 1597341371
transform 1 0 15916 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1597341371
transform 1 0 16008 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1597341371
transform 1 0 16192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1597341371
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1597341371
transform 1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _182_
timestamp 1597341371
transform 1 0 16560 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_170
timestamp 1597341371
transform 1 0 16744 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1597341371
transform 1 0 17388 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1597341371
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_177
timestamp 1597341371
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_174
timestamp 1597341371
transform 1 0 17112 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1597341371
transform 1 0 17204 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1597341371
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A2
timestamp 1597341371
transform 1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1597341371
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_183
timestamp 1597341371
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1597341371
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1597341371
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1597341371
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1597341371
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _184_
timestamp 1597341371
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_196
timestamp 1597341371
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_192
timestamp 1597341371
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1597341371
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_192
timestamp 1597341371
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__B1
timestamp 1597341371
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__B1
timestamp 1597341371
transform 1 0 18584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__B1
timestamp 1597341371
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A2
timestamp 1597341371
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__B2
timestamp 1597341371
transform 1 0 19320 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _222_
timestamp 1597341371
transform 1 0 19320 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 1597341371
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_204
timestamp 1597341371
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1597341371
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_209
timestamp 1597341371
transform 1 0 20332 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1597341371
transform 1 0 19964 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 1597341371
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__C
timestamp 1597341371
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A1
timestamp 1597341371
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A3
timestamp 1597341371
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1597341371
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1597341371
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1597341371
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1597341371
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B1
timestamp 1597341371
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1597341371
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _218_
timestamp 1597341371
transform 1 0 21160 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _226_
timestamp 1597341371
transform 1 0 21068 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_10_243
timestamp 1597341371
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_231
timestamp 1597341371
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1597341371
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1597341371
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_231
timestamp 1597341371
transform 1 0 22356 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_227
timestamp 1597341371
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__B2
timestamp 1597341371
transform 1 0 22172 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1597341371
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1597341371
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_255
timestamp 1597341371
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1597341371
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1597341371
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_292
timestamp 1597341371
transform 1 0 27968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_288
timestamp 1597341371
transform 1 0 27600 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1597341371
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1597341371
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1597341371
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1597341371
transform -1 0 28336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1597341371
transform -1 0 28336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1597341371
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1597341371
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1597341371
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1597341371
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1597341371
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1597341371
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1597341371
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1597341371
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1597341371
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1597341371
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1597341371
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1597341371
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_39
timestamp 1597341371
transform 1 0 4692 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1597341371
transform 1 0 5152 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__B1
timestamp 1597341371
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1597341371
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1597341371
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1597341371
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1597341371
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1597341371
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1597341371
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_51
timestamp 1597341371
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1597341371
transform 1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1597341371
transform 1 0 5980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1597341371
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1597341371
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1597341371
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 1597341371
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A1
timestamp 1597341371
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1597341371
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1597341371
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1597341371
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1597341371
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__RESET_B
timestamp 1597341371
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1597341371
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1597341371
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1597341371
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1597341371
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _142_
timestamp 1597341371
transform 1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_73
timestamp 1597341371
transform 1 0 7820 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_69
timestamp 1597341371
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1597341371
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 1597341371
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__B2
timestamp 1597341371
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__D
timestamp 1597341371
transform 1 0 7636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__CLK
timestamp 1597341371
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _186_
timestamp 1597341371
transform 1 0 7084 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_4  _295_
timestamp 1597341371
transform 1 0 6992 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_12_84
timestamp 1597341371
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_76
timestamp 1597341371
transform 1 0 8096 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _192_
timestamp 1597341371
transform 1 0 8188 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1597341371
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1597341371
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1597341371
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1597341371
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1597341371
transform 1 0 9568 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A2
timestamp 1597341371
transform 1 0 9292 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B2
timestamp 1597341371
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__CLK
timestamp 1597341371
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1597341371
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1597341371
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1597341371
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_96
timestamp 1597341371
transform 1 0 9936 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B1
timestamp 1597341371
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _172_
timestamp 1597341371
transform 1 0 9844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _193_
timestamp 1597341371
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _190_
timestamp 1597341371
transform 1 0 10028 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1597341371
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1597341371
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1597341371
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A1
timestamp 1597341371
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__D
timestamp 1597341371
transform 1 0 10672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _185_
timestamp 1597341371
transform 1 0 10764 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _170_
timestamp 1597341371
transform 1 0 11040 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1597341371
transform 1 0 11960 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1597341371
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_119
timestamp 1597341371
transform 1 0 12052 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1597341371
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1597341371
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1597341371
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A3
timestamp 1597341371
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B
timestamp 1597341371
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__RESET_B
timestamp 1597341371
transform 1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1597341371
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1597341371
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1597341371
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1597341371
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1597341371
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1597341371
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1597341371
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1597341371
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A2
timestamp 1597341371
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A1
timestamp 1597341371
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1597341371
transform 1 0 13340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1597341371
transform 1 0 14536 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_145
timestamp 1597341371
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1597341371
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1597341371
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B1
timestamp 1597341371
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _261_
timestamp 1597341371
transform 1 0 13708 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _296_
timestamp 1597341371
transform 1 0 12880 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__o21a_4  _266_
timestamp 1597341371
transform 1 0 12972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1597341371
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1597341371
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1597341371
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_151
timestamp 1597341371
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1597341371
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1597341371
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__B
timestamp 1597341371
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1597341371
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_156
timestamp 1597341371
transform 1 0 15456 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_161
timestamp 1597341371
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1597341371
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1597341371
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__B2
timestamp 1597341371
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _209_
timestamp 1597341371
transform 1 0 15732 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_169
timestamp 1597341371
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1597341371
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1597341371
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_168
timestamp 1597341371
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1_N
timestamp 1597341371
transform 1 0 16468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A2_N
timestamp 1597341371
transform 1 0 16100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__CLK
timestamp 1597341371
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _280_
timestamp 1597341371
transform 1 0 16836 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__a2bb2o_4  _267_
timestamp 1597341371
transform 1 0 15732 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_175
timestamp 1597341371
transform 1 0 17204 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1597341371
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__D
timestamp 1597341371
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1597341371
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1597341371
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1597341371
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__RESET_B
timestamp 1597341371
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1597341371
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1597341371
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1597341371
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1597341371
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _198_
timestamp 1597341371
transform 1 0 18216 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_198
timestamp 1597341371
transform 1 0 19320 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1597341371
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1597341371
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_193
timestamp 1597341371
transform 1 0 18860 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1597341371
transform 1 0 18492 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1597341371
transform 1 0 18952 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__D
timestamp 1597341371
transform 1 0 19136 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _220_
timestamp 1597341371
transform 1 0 18400 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_4  _212_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 19320 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_13_204
timestamp 1597341371
transform 1 0 19872 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1597341371
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1597341371
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_205
timestamp 1597341371
transform 1 0 19964 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1597341371
transform 1 0 19688 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1597341371
transform 1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _225_
timestamp 1597341371
transform 1 0 20240 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _217_
timestamp 1597341371
transform 1 0 19688 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_223
timestamp 1597341371
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_217
timestamp 1597341371
transform 1 0 21068 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1597341371
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_220
timestamp 1597341371
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1597341371
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__B2
timestamp 1597341371
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__B
timestamp 1597341371
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__RESET_B
timestamp 1597341371
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1597341371
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _227_
timestamp 1597341371
transform 1 0 21068 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_224
timestamp 1597341371
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1_N
timestamp 1597341371
transform 1 0 21896 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _157_
timestamp 1597341371
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1597341371
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_228
timestamp 1597341371
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A2_N
timestamp 1597341371
transform 1 0 22264 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__CLK
timestamp 1597341371
transform 1 0 22264 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_232
timestamp 1597341371
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_233
timestamp 1597341371
transform 1 0 22540 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_232
timestamp 1597341371
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__B1
timestamp 1597341371
transform 1 0 22632 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1597341371
transform 1 0 22724 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__D
timestamp 1597341371
transform 1 0 22632 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1597341371
transform 1 0 23184 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1597341371
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_237
timestamp 1597341371
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_236
timestamp 1597341371
transform 1 0 22816 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A2
timestamp 1597341371
transform 1 0 23000 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__D
timestamp 1597341371
transform 1 0 23092 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1597341371
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1597341371
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1597341371
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_241
timestamp 1597341371
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1597341371
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1597341371
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1597341371
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1597341371
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_265
timestamp 1597341371
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1597341371
transform 1 0 24380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1597341371
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1597341371
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1597341371
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_292
timestamp 1597341371
transform 1 0 27968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_288
timestamp 1597341371
transform 1 0 27600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1597341371
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1597341371
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1597341371
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1597341371
transform -1 0 28336 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1597341371
transform -1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1597341371
transform -1 0 28336 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1597341371
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1597341371
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1597341371
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1597341371
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1597341371
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1597341371
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1597341371
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1597341371
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_44
timestamp 1597341371
transform 1 0 5152 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1597341371
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1597341371
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1597341371
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1597341371
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1597341371
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1597341371
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1597341371
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_52
timestamp 1597341371
transform 1 0 5888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1597341371
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A3
timestamp 1597341371
transform 1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1597341371
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _188_
timestamp 1597341371
transform 1 0 6164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1597341371
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_66
timestamp 1597341371
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1597341371
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__B2
timestamp 1597341371
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1597341371
transform 1 0 6992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A2_N
timestamp 1597341371
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _194_
timestamp 1597341371
transform 1 0 7176 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1597341371
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_83
timestamp 1597341371
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A1_N
timestamp 1597341371
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_97
timestamp 1597341371
transform 1 0 10028 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1597341371
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_99
timestamp 1597341371
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1597341371
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1597341371
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1597341371
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__B1
timestamp 1597341371
transform 1 0 9844 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1597341371
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1597341371
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _189_
timestamp 1597341371
transform 1 0 8188 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_109
timestamp 1597341371
transform 1 0 11132 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_105
timestamp 1597341371
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_101
timestamp 1597341371
transform 1 0 10396 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1597341371
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1597341371
transform 1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1597341371
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1597341371
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_124
timestamp 1597341371
transform 1 0 12512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1597341371
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1597341371
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _294_
timestamp 1597341371
transform 1 0 10396 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_15_127
timestamp 1597341371
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_128
timestamp 1597341371
transform 1 0 12880 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1597341371
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1597341371
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B2
timestamp 1597341371
transform 1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__B1
timestamp 1597341371
transform 1 0 13064 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1597341371
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_135
timestamp 1597341371
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A1
timestamp 1597341371
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__RESET_B
timestamp 1597341371
transform 1 0 13340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1597341371
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1597341371
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1597341371
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1597341371
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__D
timestamp 1597341371
transform 1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__CLK
timestamp 1597341371
transform 1 0 14168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp 1597341371
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _288_
timestamp 1597341371
transform 1 0 13800 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1597341371
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1597341371
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1597341371
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _183_
timestamp 1597341371
transform 1 0 15456 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1597341371
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1597341371
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1597341371
transform 1 0 16100 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1597341371
transform 1 0 16652 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_165
timestamp 1597341371
transform 1 0 16284 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1597341371
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1597341371
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _246_
timestamp 1597341371
transform 1 0 16652 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _224_
timestamp 1597341371
transform 1 0 16744 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1597341371
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1597341371
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1597341371
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_180
timestamp 1597341371
transform 1 0 17664 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_176
timestamp 1597341371
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__C
timestamp 1597341371
transform 1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B
timestamp 1597341371
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__B
timestamp 1597341371
transform 1 0 17940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A1
timestamp 1597341371
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1597341371
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1597341371
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1597341371
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 1597341371
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__C
timestamp 1597341371
transform 1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _219_
timestamp 1597341371
transform 1 0 18676 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _210_
timestamp 1597341371
transform 1 0 18216 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_195
timestamp 1597341371
transform 1 0 19044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__B
timestamp 1597341371
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_204
timestamp 1597341371
transform 1 0 19872 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1597341371
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1597341371
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_204
timestamp 1597341371
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_200
timestamp 1597341371
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__B
timestamp 1597341371
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A
timestamp 1597341371
transform 1 0 19688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__B1
timestamp 1597341371
transform 1 0 20240 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1597341371
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1597341371
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_219
timestamp 1597341371
transform 1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1597341371
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__D
timestamp 1597341371
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__C1
timestamp 1597341371
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1597341371
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _257_
timestamp 1597341371
transform 1 0 20240 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_15_234
timestamp 1597341371
transform 1 0 22632 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1597341371
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_226
timestamp 1597341371
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A1
timestamp 1597341371
transform 1 0 22080 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A2
timestamp 1597341371
transform 1 0 21712 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1597341371
transform 1 0 22448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_238
timestamp 1597341371
transform 1 0 23000 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1597341371
transform 1 0 22816 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1597341371
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1597341371
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_248
timestamp 1597341371
transform 1 0 23920 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _283_
timestamp 1597341371
transform 1 0 21804 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1597341371
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1597341371
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_272
timestamp 1597341371
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_260
timestamp 1597341371
transform 1 0 25024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1597341371
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_292
timestamp 1597341371
transform 1 0 27968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_288
timestamp 1597341371
transform 1 0 27600 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1597341371
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1597341371
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1597341371
transform -1 0 28336 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1597341371
transform -1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1597341371
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1597341371
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1597341371
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1597341371
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1597341371
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1597341371
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1597341371
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1597341371
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1597341371
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1597341371
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1597341371
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1597341371
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1597341371
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1597341371
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_56
timestamp 1597341371
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1597341371
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _191_
timestamp 1597341371
transform 1 0 6440 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1597341371
transform 1 0 7912 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1597341371
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1597341371
transform 1 0 7268 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1597341371
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1597341371
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_94
timestamp 1597341371
transform 1 0 9752 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1597341371
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1597341371
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1597341371
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1597341371
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__B
timestamp 1597341371
transform 1 0 9016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1597341371
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _187_
timestamp 1597341371
transform 1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _176_
timestamp 1597341371
transform 1 0 8004 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1597341371
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A2
timestamp 1597341371
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1597341371
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1597341371
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1597341371
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__CLK
timestamp 1597341371
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp 1597341371
transform 1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1597341371
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__B1
timestamp 1597341371
transform 1 0 11500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__D
timestamp 1597341371
transform 1 0 11408 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1597341371
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1597341371
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_115
timestamp 1597341371
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__RESET_B
timestamp 1597341371
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _164_
timestamp 1597341371
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1597341371
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_120
timestamp 1597341371
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A1
timestamp 1597341371
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1597341371
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_133
timestamp 1597341371
transform 1 0 13340 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1597341371
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1597341371
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__B1
timestamp 1597341371
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__B2
timestamp 1597341371
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A3
timestamp 1597341371
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1597341371
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1597341371
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1597341371
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1597341371
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1597341371
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__C1
timestamp 1597341371
transform 1 0 13984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A2
timestamp 1597341371
transform 1 0 14352 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__B1_N
timestamp 1597341371
transform 1 0 14352 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A1
timestamp 1597341371
transform 1 0 14720 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _256_
timestamp 1597341371
transform 1 0 14720 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_4  _251_
timestamp 1597341371
transform 1 0 12604 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1597341371
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1597341371
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1597341371
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A3
timestamp 1597341371
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1597341371
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _211_
timestamp 1597341371
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1597341371
transform 1 0 16652 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 1597341371
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1597341371
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__C
timestamp 1597341371
transform 1 0 16468 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A2
timestamp 1597341371
transform 1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _252_
timestamp 1597341371
transform 1 0 16468 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1597341371
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1597341371
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1597341371
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1597341371
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1597341371
transform 1 0 17572 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A2_N
timestamp 1597341371
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B1
timestamp 1597341371
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1597341371
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_189
timestamp 1597341371
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_193
timestamp 1597341371
transform 1 0 18860 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1597341371
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1597341371
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1_N
timestamp 1597341371
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__B1
timestamp 1597341371
transform 1 0 18676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _263_
timestamp 1597341371
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _258_
timestamp 1597341371
transform 1 0 18676 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_211
timestamp 1597341371
transform 1 0 20516 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_207
timestamp 1597341371
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1597341371
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A
timestamp 1597341371
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A1
timestamp 1597341371
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1597341371
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1597341371
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1597341371
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _229_
timestamp 1597341371
transform 1 0 21068 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _260_
timestamp 1597341371
transform 1 0 20884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_235
timestamp 1597341371
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1597341371
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_227
timestamp 1597341371
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_230
timestamp 1597341371
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_226
timestamp 1597341371
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__B
timestamp 1597341371
transform 1 0 22540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 1597341371
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__B1
timestamp 1597341371
transform 1 0 22080 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _259_
timestamp 1597341371
transform 1 0 22448 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1597341371
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1597341371
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1597341371
transform 1 0 23092 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A1
timestamp 1597341371
transform 1 0 22908 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1597341371
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_241
timestamp 1597341371
transform 1 0 23276 0 -1 11424
box -38 -48 1142 592
use AMUX2_3V  AMUX2_3V
timestamp 1598931070
transform 1 0 23828 0 1 11424
box 0 -48 1748 1136
use sky130_fd_sc_hd__decap_12  FILLER_17_266
timestamp 1597341371
transform 1 0 25576 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_273
timestamp 1597341371
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_265
timestamp 1597341371
transform 1 0 25484 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1597341371
transform 1 0 24380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_290
timestamp 1597341371
transform 1 0 27784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_278
timestamp 1597341371
transform 1 0 26680 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_292
timestamp 1597341371
transform 1 0 27968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_288
timestamp 1597341371
transform 1 0 27600 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1597341371
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1597341371
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1597341371
transform -1 0 28336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1597341371
transform -1 0 28336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1597341371
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1597341371
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1597341371
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1597341371
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1597341371
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1597341371
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1597341371
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1597341371
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1597341371
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1597341371
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1597341371
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1597341371
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1597341371
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1597341371
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1597341371
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1597341371
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1597341371
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1597341371
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1597341371
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1597341371
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1597341371
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_93
timestamp 1597341371
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1597341371
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1597341371
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1597341371
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_101
timestamp 1597341371
transform 1 0 10396 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A1
timestamp 1597341371
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__B
timestamp 1597341371
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1597341371
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1597341371
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1597341371
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1597341371
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A1
timestamp 1597341371
transform 1 0 11592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__B1
timestamp 1597341371
transform 1 0 11960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1597341371
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _287_
timestamp 1597341371
transform 1 0 11040 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1597341371
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1597341371
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__B1
timestamp 1597341371
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_143
timestamp 1597341371
transform 1 0 14260 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1597341371
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1597341371
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_143
timestamp 1597341371
transform 1 0 14260 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_139
timestamp 1597341371
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A2
timestamp 1597341371
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A2
timestamp 1597341371
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A1
timestamp 1597341371
transform 1 0 13708 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__B1
timestamp 1597341371
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _255_
timestamp 1597341371
transform 1 0 14628 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ai_4  _250_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 12696 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1597341371
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1597341371
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1597341371
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1597341371
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1597341371
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_165
timestamp 1597341371
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1597341371
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A2
timestamp 1597341371
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__B
timestamp 1597341371
transform 1 0 16468 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__B1
timestamp 1597341371
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__B
timestamp 1597341371
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__a21boi_4  _254_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 15456 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1597341371
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1597341371
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1597341371
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1597341371
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__D
timestamp 1597341371
transform 1 0 17204 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B1
timestamp 1597341371
transform 1 0 17572 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1597341371
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1597341371
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_194
timestamp 1597341371
transform 1 0 18952 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1597341371
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__C
timestamp 1597341371
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A1
timestamp 1597341371
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _238_
timestamp 1597341371
transform 1 0 19320 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _231_
timestamp 1597341371
transform 1 0 18768 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _248_
timestamp 1597341371
transform 1 0 17388 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1597341371
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 1597341371
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1597341371
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A2
timestamp 1597341371
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 1597341371
transform 1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B2
timestamp 1597341371
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1597341371
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1597341371
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1597341371
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1597341371
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__B2
timestamp 1597341371
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1597341371
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1597341371
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 1597341371
transform 1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A2
timestamp 1597341371
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1597341371
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1597341371
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_219
timestamp 1597341371
transform 1 0 21252 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__RESET_B
timestamp 1597341371
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _264_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 21436 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1597341371
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_230
timestamp 1597341371
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__D
timestamp 1597341371
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1597341371
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1597341371
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_238
timestamp 1597341371
transform 1 0 23000 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__B1
timestamp 1597341371
transform 1 0 22816 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__CLK
timestamp 1597341371
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1597341371
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_245
timestamp 1597341371
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_242
timestamp 1597341371
transform 1 0 23368 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_AMUX2_3V_select
timestamp 1597341371
transform 1 0 23460 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1597341371
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_AMUX2_3V_I1
timestamp 1597341371
transform 1 0 23828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _265_
timestamp 1597341371
transform 1 0 21712 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_273
timestamp 1597341371
transform 1 0 26220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1597341371
transform 1 0 25116 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1597341371
transform 1 0 24012 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_266
timestamp 1597341371
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_285
timestamp 1597341371
transform 1 0 27324 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_292
timestamp 1597341371
transform 1 0 27968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1597341371
transform 1 0 27600 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1597341371
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1597341371
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1597341371
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1597341371
transform -1 0 28336 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1597341371
transform -1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1597341371
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1597341371
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1597341371
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1597341371
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1597341371
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1597341371
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1597341371
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1597341371
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1597341371
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1597341371
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1597341371
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1597341371
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_74
timestamp 1597341371
transform 1 0 7912 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1597341371
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1597341371
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1597341371
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1597341371
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1597341371
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1597341371
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_80
timestamp 1597341371
transform 1 0 8464 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_83
timestamp 1597341371
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1597341371
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1597341371
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _175_
timestamp 1597341371
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1597341371
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1597341371
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_96
timestamp 1597341371
transform 1 0 9936 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_84
timestamp 1597341371
transform 1 0 8832 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1597341371
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_108
timestamp 1597341371
transform 1 0 11040 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_107
timestamp 1597341371
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B1
timestamp 1597341371
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A2
timestamp 1597341371
transform 1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B2
timestamp 1597341371
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_111
timestamp 1597341371
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp 1597341371
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A3
timestamp 1597341371
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__D
timestamp 1597341371
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1597341371
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1597341371
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__RESET_B
timestamp 1597341371
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__CLK
timestamp 1597341371
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1597341371
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1597341371
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1597341371
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 1597341371
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1597341371
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_125
timestamp 1597341371
transform 1 0 12604 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_147
timestamp 1597341371
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_142
timestamp 1597341371
transform 1 0 14168 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1597341371
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_144
timestamp 1597341371
transform 1 0 14352 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_140
timestamp 1597341371
transform 1 0 13984 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1597341371
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A
timestamp 1597341371
transform 1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__C
timestamp 1597341371
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _253_
timestamp 1597341371
transform 1 0 14812 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _247_
timestamp 1597341371
transform 1 0 12604 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_4  _245_
timestamp 1597341371
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1597341371
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1597341371
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1597341371
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1597341371
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _262_
timestamp 1597341371
transform 1 0 15456 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_162
timestamp 1597341371
transform 1 0 16008 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_165
timestamp 1597341371
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A
timestamp 1597341371
transform 1 0 16468 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1597341371
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _239_
timestamp 1597341371
transform 1 0 16376 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1597341371
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _249_ home/praharsha/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597341371
transform 1 0 16836 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1597341371
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1597341371
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1597341371
transform 1 0 17204 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1597341371
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1597341371
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A2
timestamp 1597341371
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B2
timestamp 1597341371
transform 1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B1
timestamp 1597341371
transform 1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1597341371
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1597341371
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _234_
timestamp 1597341371
transform 1 0 18400 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _230_
timestamp 1597341371
transform 1 0 18584 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1597341371
transform 1 0 20056 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1597341371
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp 1597341371
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1597341371
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1597341371
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 1597341371
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1597341371
transform 1 0 19872 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _232_
timestamp 1597341371
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1597341371
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1597341371
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1597341371
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__D
timestamp 1597341371
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1597341371
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1597341371
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1597341371
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__C
timestamp 1597341371
transform 1 0 21068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1597341371
transform 1 0 21252 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_223
timestamp 1597341371
transform 1 0 21620 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_221
timestamp 1597341371
transform 1 0 21436 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1597341371
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_241
timestamp 1597341371
transform 1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_233
timestamp 1597341371
transform 1 0 22540 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_226
timestamp 1597341371
transform 1 0 21896 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A1
timestamp 1597341371
transform 1 0 21712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1597341371
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _297_
timestamp 1597341371
transform 1 0 22264 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1597341371
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1597341371
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_273
timestamp 1597341371
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_265
timestamp 1597341371
transform 1 0 25484 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1597341371
transform 1 0 24380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1597341371
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_292
timestamp 1597341371
transform 1 0 27968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_288
timestamp 1597341371
transform 1 0 27600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1597341371
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1597341371
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1597341371
transform -1 0 28336 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1597341371
transform -1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1597341371
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1597341371
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1597341371
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1597341371
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1597341371
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1597341371
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1597341371
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1597341371
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1597341371
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1597341371
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1597341371
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1597341371
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1597341371
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1597341371
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1597341371
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1597341371
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1597341371
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1597341371
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1597341371
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1597341371
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1597341371
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1597341371
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1597341371
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1597341371
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1597341371
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1597341371
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1597341371
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1597341371
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _286_
timestamp 1597341371
transform 1 0 11868 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_23_128
timestamp 1597341371
transform 1 0 12880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1597341371
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _244_
timestamp 1597341371
transform 1 0 13156 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_140
timestamp 1597341371
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_140
timestamp 1597341371
transform 1 0 13984 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1597341371
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1597341371
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1597341371
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1597341371
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_144
timestamp 1597341371
transform 1 0 14352 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A
timestamp 1597341371
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1597341371
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B
timestamp 1597341371
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1597341371
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1597341371
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1597341371
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1597341371
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _236_
timestamp 1597341371
transform 1 0 14904 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1597341371
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_163
timestamp 1597341371
transform 1 0 16100 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1597341371
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__B
timestamp 1597341371
transform 1 0 17020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A2
timestamp 1597341371
transform 1 0 16192 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _240_
timestamp 1597341371
transform 1 0 16560 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _243_
timestamp 1597341371
transform 1 0 15640 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1597341371
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1597341371
transform 1 0 17204 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1597341371
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1597341371
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1597341371
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_179
timestamp 1597341371
transform 1 0 17572 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A2_N
timestamp 1597341371
transform 1 0 17848 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1597341371
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1597341371
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1597341371
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1_N
timestamp 1597341371
transform 1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_190
timestamp 1597341371
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1597341371
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A
timestamp 1597341371
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _228_
timestamp 1597341371
transform 1 0 18768 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _235_
timestamp 1597341371
transform 1 0 18584 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1597341371
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_201
timestamp 1597341371
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1597341371
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_206
timestamp 1597341371
transform 1 0 20056 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B2
timestamp 1597341371
transform 1 0 19780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__CLK
timestamp 1597341371
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1597341371
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_215
timestamp 1597341371
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__RESET_B
timestamp 1597341371
transform 1 0 21620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1597341371
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1597341371
transform 1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _284_
timestamp 1597341371
transform 1 0 20332 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1597341371
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1597341371
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1597341371
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1597341371
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1597341371
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1597341371
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1597341371
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_273
timestamp 1597341371
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_261
timestamp 1597341371
transform 1 0 25116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_249
timestamp 1597341371
transform 1 0 24012 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1597341371
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_292
timestamp 1597341371
transform 1 0 27968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_288
timestamp 1597341371
transform 1 0 27600 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1597341371
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1597341371
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1597341371
transform -1 0 28336 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1597341371
transform -1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1597341371
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1597341371
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1597341371
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1597341371
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1597341371
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1597341371
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1597341371
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1597341371
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1597341371
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1597341371
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1597341371
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1597341371
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1597341371
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1597341371
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1597341371
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1597341371
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1597341371
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1597341371
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1597341371
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1597341371
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1597341371
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1597341371
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1597341371
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1597341371
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1597341371
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1597341371
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1597341371
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1597341371
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1597341371
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1597341371
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1597341371
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1597341371
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1597341371
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1597341371
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1597341371
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1597341371
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1597341371
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1597341371
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1597341371
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1597341371
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_117
timestamp 1597341371
transform 1 0 11868 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1597341371
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1597341371
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_135
timestamp 1597341371
transform 1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_133
timestamp 1597341371
transform 1 0 13340 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1597341371
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_125
timestamp 1597341371
transform 1 0 12604 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1597341371
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _154_
timestamp 1597341371
transform 1 0 12696 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_140
timestamp 1597341371
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1597341371
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_137
timestamp 1597341371
transform 1 0 13708 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1597341371
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__RESET_B
timestamp 1597341371
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__CLK
timestamp 1597341371
transform 1 0 14168 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1597341371
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1597341371
transform 1 0 14720 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1597341371
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__D
timestamp 1597341371
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_144
timestamp 1597341371
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1597341371
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _285_
timestamp 1597341371
transform 1 0 14168 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1597341371
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1597341371
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1597341371
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1597341371
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1597341371
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1597341371
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _242_
timestamp 1597341371
transform 1 0 15456 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _237_
timestamp 1597341371
transform 1 0 15456 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_25_173
timestamp 1597341371
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1597341371
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1597341371
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1597341371
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_163
timestamp 1597341371
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B1
timestamp 1597341371
transform 1 0 16376 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__B
timestamp 1597341371
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__A
timestamp 1597341371
transform 1 0 16468 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_163
timestamp 1597341371
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _241_
timestamp 1597341371
transform 1 0 16744 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 1597341371
transform 1 0 17388 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1597341371
transform 1 0 18032 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__B2
timestamp 1597341371
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1597341371
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1597341371
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1597341371
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _233_
timestamp 1597341371
transform 1 0 18768 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_187
timestamp 1597341371
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_175
timestamp 1597341371
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1597341371
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1597341371
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1597341371
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1597341371
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1597341371
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1597341371
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1597341371
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_199
timestamp 1597341371
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1597341371
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1597341371
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1597341371
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1597341371
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1597341371
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1597341371
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1597341371
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1597341371
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1597341371
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1597341371
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1597341371
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1597341371
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1597341371
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1597341371
transform 1 0 25852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1597341371
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1597341371
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1597341371
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1597341371
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1597341371
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_292
timestamp 1597341371
transform 1 0 27968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1597341371
transform 1 0 27600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1597341371
transform 1 0 27968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_288
timestamp 1597341371
transform 1 0 27600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1597341371
transform -1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1597341371
transform -1 0 28336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1597341371
transform -1 0 28336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1597341371
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1597341371
transform 1 0 26956 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1597341371
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1597341371
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1597341371
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1597341371
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1597341371
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1597341371
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1597341371
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1597341371
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1597341371
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1597341371
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1597341371
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1597341371
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1597341371
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1597341371
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1597341371
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1597341371
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1597341371
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1597341371
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1597341371
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1597341371
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1597341371
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1597341371
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1597341371
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1597341371
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1597341371
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1597341371
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1597341371
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1597341371
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1597341371
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1597341371
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1597341371
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1597341371
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1597341371
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1597341371
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1597341371
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1597341371
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1597341371
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1597341371
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1597341371
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1597341371
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1597341371
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1597341371
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1597341371
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1597341371
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1597341371
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1597341371
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1597341371
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1597341371
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1597341371
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1597341371
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1597341371
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1597341371
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1597341371
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1597341371
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1597341371
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1597341371
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1597341371
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1597341371
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_292
timestamp 1597341371
transform 1 0 27968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1597341371
transform 1 0 27600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1597341371
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1597341371
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1597341371
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1597341371
transform -1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1597341371
transform -1 0 28336 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1597341371
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1597341371
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1597341371
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1597341371
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1597341371
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1597341371
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1597341371
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1597341371
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1597341371
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1597341371
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1597341371
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1597341371
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1597341371
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1597341371
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1597341371
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1597341371
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1597341371
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1597341371
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1597341371
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1597341371
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1597341371
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1597341371
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1597341371
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1597341371
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1597341371
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1597341371
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1597341371
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1597341371
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1597341371
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1597341371
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1597341371
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1597341371
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1597341371
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1597341371
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1597341371
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1597341371
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1597341371
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1597341371
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1597341371
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1597341371
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1597341371
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1597341371
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1597341371
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1597341371
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1597341371
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1597341371
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1597341371
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1597341371
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1597341371
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1597341371
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1597341371
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1597341371
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1597341371
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1597341371
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1597341371
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1597341371
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1597341371
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_292
timestamp 1597341371
transform 1 0 27968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_288
timestamp 1597341371
transform 1 0 27600 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1597341371
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1597341371
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1597341371
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1597341371
transform -1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1597341371
transform -1 0 28336 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1597341371
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1597341371
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1597341371
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1597341371
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1597341371
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1597341371
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1597341371
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1597341371
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1597341371
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1597341371
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1597341371
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1597341371
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1597341371
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1597341371
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1597341371
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1597341371
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1597341371
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1597341371
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1597341371
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1597341371
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1597341371
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1597341371
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1597341371
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1597341371
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1597341371
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1597341371
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1597341371
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1597341371
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1597341371
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1597341371
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1597341371
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1597341371
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1597341371
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1597341371
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1597341371
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1597341371
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1597341371
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1597341371
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1597341371
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1597341371
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1597341371
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1597341371
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1597341371
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1597341371
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1597341371
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1597341371
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1597341371
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1597341371
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1597341371
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1597341371
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1597341371
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1597341371
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1597341371
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1597341371
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1597341371
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1597341371
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1597341371
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_292
timestamp 1597341371
transform 1 0 27968 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1597341371
transform 1 0 27600 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1597341371
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1597341371
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1597341371
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1597341371
transform -1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1597341371
transform -1 0 28336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1597341371
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1597341371
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1597341371
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1597341371
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1597341371
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1597341371
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1597341371
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1597341371
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1597341371
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1597341371
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1597341371
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1597341371
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1597341371
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1597341371
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1597341371
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1597341371
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1597341371
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1597341371
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1597341371
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1597341371
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1597341371
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1597341371
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1597341371
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1597341371
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1597341371
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1597341371
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1597341371
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1597341371
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1597341371
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1597341371
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1597341371
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1597341371
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1597341371
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1597341371
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1597341371
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1597341371
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1597341371
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1597341371
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1597341371
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1597341371
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1597341371
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1597341371
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1597341371
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1597341371
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1597341371
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1597341371
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1597341371
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1597341371
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1597341371
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1597341371
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1597341371
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1597341371
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1597341371
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1597341371
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1597341371
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1597341371
transform 1 0 25852 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1597341371
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_292
timestamp 1597341371
transform 1 0 27968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1597341371
transform 1 0 27600 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1597341371
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1597341371
transform 1 0 26956 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1597341371
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1597341371
transform -1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1597341371
transform -1 0 28336 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1597341371
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1597341371
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1597341371
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1597341371
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1597341371
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1597341371
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1597341371
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1597341371
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1597341371
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1597341371
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1597341371
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1597341371
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1597341371
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1597341371
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1597341371
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1597341371
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1597341371
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1597341371
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1597341371
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1597341371
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1597341371
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1597341371
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1597341371
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1597341371
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1597341371
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1597341371
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1597341371
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1597341371
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1597341371
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1597341371
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1597341371
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1597341371
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1597341371
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1597341371
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1597341371
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1597341371
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1597341371
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1597341371
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1597341371
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1597341371
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1597341371
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1597341371
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1597341371
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1597341371
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1597341371
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1597341371
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1597341371
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1597341371
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1597341371
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1597341371
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1597341371
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1597341371
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1597341371
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1597341371
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1597341371
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1597341371
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1597341371
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1597341371
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1597341371
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1597341371
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1597341371
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1597341371
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1597341371
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1597341371
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1597341371
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1597341371
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1597341371
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1597341371
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1597341371
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1597341371
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1597341371
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1597341371
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1597341371
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1597341371
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1597341371
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1597341371
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1597341371
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1597341371
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1597341371
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1597341371
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_269
timestamp 1597341371
transform 1 0 25852 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1597341371
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1597341371
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1597341371
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_269
timestamp 1597341371
transform 1 0 25852 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1597341371
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1597341371
transform 1 0 26956 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_292
timestamp 1597341371
transform 1 0 27968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1597341371
transform 1 0 27600 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1597341371
transform 1 0 26496 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1597341371
transform 1 0 26956 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1597341371
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1597341371
transform -1 0 28336 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1597341371
transform -1 0 28336 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1597341371
transform -1 0 28336 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1597341371
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1597341371
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1597341371
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1597341371
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1597341371
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1597341371
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1597341371
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1597341371
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1597341371
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1597341371
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1597341371
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1597341371
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1597341371
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1597341371
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1597341371
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1597341371
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1597341371
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1597341371
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1597341371
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1597341371
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1597341371
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1597341371
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1597341371
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1597341371
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1597341371
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1597341371
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1597341371
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1597341371
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1597341371
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1597341371
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1597341371
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1597341371
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1597341371
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1597341371
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1597341371
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1597341371
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1597341371
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1597341371
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1597341371
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1597341371
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1597341371
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1597341371
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1597341371
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1597341371
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1597341371
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1597341371
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1597341371
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1597341371
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1597341371
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1597341371
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1597341371
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1597341371
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1597341371
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1597341371
transform 1 0 25852 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1597341371
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1597341371
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1597341371
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1597341371
transform 1 0 26956 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_292
timestamp 1597341371
transform 1 0 27968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1597341371
transform 1 0 27600 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1597341371
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1597341371
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1597341371
transform -1 0 28336 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1597341371
transform -1 0 28336 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1597341371
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1597341371
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1597341371
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1597341371
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1597341371
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1597341371
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1597341371
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1597341371
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1597341371
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1597341371
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1597341371
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1597341371
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1597341371
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1597341371
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1597341371
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1597341371
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1597341371
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1597341371
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1597341371
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1597341371
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1597341371
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1597341371
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1597341371
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1597341371
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1597341371
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1597341371
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1597341371
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1597341371
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1597341371
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1597341371
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1597341371
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1597341371
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1597341371
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1597341371
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1597341371
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1597341371
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1597341371
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1597341371
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1597341371
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1597341371
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1597341371
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1597341371
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1597341371
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1597341371
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1597341371
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1597341371
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1597341371
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1597341371
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1597341371
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1597341371
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1597341371
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1597341371
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1597341371
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_269
timestamp 1597341371
transform 1 0 25852 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1597341371
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1597341371
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1597341371
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1597341371
transform 1 0 26956 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_292
timestamp 1597341371
transform 1 0 27968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1597341371
transform 1 0 27600 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1597341371
transform 1 0 26496 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1597341371
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1597341371
transform -1 0 28336 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1597341371
transform -1 0 28336 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1597341371
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1597341371
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1597341371
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1597341371
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1597341371
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1597341371
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1597341371
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1597341371
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1597341371
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1597341371
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1597341371
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1597341371
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_74
timestamp 1597341371
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1597341371
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1597341371
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_51
timestamp 1597341371
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1597341371
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1597341371
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1597341371
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_98
timestamp 1597341371
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_86
timestamp 1597341371
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1597341371
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_80
timestamp 1597341371
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1597341371
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1597341371
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_110
timestamp 1597341371
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_117
timestamp 1597341371
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1597341371
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1597341371
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_147
timestamp 1597341371
transform 1 0 14628 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1597341371
transform 1 0 13524 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1597341371
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1597341371
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_171
timestamp 1597341371
transform 1 0 16836 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_159
timestamp 1597341371
transform 1 0 15732 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_166
timestamp 1597341371
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1597341371
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1597341371
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1597341371
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1597341371
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_190
timestamp 1597341371
transform 1 0 18584 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_178
timestamp 1597341371
transform 1 0 17480 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1597341371
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1597341371
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1597341371
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1597341371
transform 1 0 20884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_202
timestamp 1597341371
transform 1 0 19688 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1597341371
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1597341371
transform 1 0 23644 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1597341371
transform 1 0 22448 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1597341371
transform 1 0 23092 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1597341371
transform 1 0 21988 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1597341371
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_269
timestamp 1597341371
transform 1 0 25852 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1597341371
transform 1 0 24748 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1597341371
transform 1 0 25300 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_251
timestamp 1597341371
transform 1 0 24196 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1597341371
transform 1 0 26956 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_292
timestamp 1597341371
transform 1 0 27968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_288
timestamp 1597341371
transform 1 0 27600 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1597341371
transform 1 0 26496 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1597341371
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1597341371
transform -1 0 28336 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1597341371
transform -1 0 28336 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1597341371
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1597341371
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1597341371
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1597341371
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1597341371
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1597341371
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1597341371
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1597341371
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1597341371
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1597341371
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1597341371
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1597341371
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_74
timestamp 1597341371
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_62
timestamp 1597341371
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1597341371
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_51
timestamp 1597341371
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1597341371
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_56
timestamp 1597341371
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1597341371
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_98
timestamp 1597341371
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_86
timestamp 1597341371
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1597341371
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_80
timestamp 1597341371
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1597341371
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1597341371
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_110
timestamp 1597341371
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1597341371
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1597341371
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1597341371
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_147
timestamp 1597341371
transform 1 0 14628 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_135
timestamp 1597341371
transform 1 0 13524 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1597341371
transform 1 0 14076 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1597341371
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1597341371
transform 1 0 16836 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_159
timestamp 1597341371
transform 1 0 15732 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_166
timestamp 1597341371
transform 1 0 16376 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1597341371
transform 1 0 15272 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1597341371
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1597341371
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1597341371
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_190
timestamp 1597341371
transform 1 0 18584 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_178
timestamp 1597341371
transform 1 0 17480 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1597341371
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_220
timestamp 1597341371
transform 1 0 21344 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1597341371
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1597341371
transform 1 0 20884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_202
timestamp 1597341371
transform 1 0 19688 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1597341371
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1597341371
transform 1 0 23644 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1597341371
transform 1 0 23184 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_232
timestamp 1597341371
transform 1 0 22448 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_239
timestamp 1597341371
transform 1 0 23092 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1597341371
transform 1 0 21988 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 1597341371
transform 1 0 23000 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1597341371
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_269
timestamp 1597341371
transform 1 0 25852 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_257
timestamp 1597341371
transform 1 0 24748 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_263
timestamp 1597341371
transform 1 0 25300 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_251
timestamp 1597341371
transform 1 0 24196 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1597341371
transform 1 0 26956 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_292
timestamp 1597341371
transform 1 0 27968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1597341371
transform 1 0 27600 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_276
timestamp 1597341371
transform 1 0 26496 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1597341371
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1597341371
transform -1 0 28336 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1597341371
transform -1 0 28336 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1597341371
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1597341371
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1597341371
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1597341371
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1597341371
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1597341371
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1597341371
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1597341371
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1597341371
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1597341371
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1597341371
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1597341371
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_74
timestamp 1597341371
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1597341371
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1597341371
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1597341371
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1597341371
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1597341371
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1597341371
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_98
timestamp 1597341371
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_86
timestamp 1597341371
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1597341371
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_80
timestamp 1597341371
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1597341371
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1597341371
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_110
timestamp 1597341371
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1597341371
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1597341371
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1597341371
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1597341371
transform 1 0 14628 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_135
timestamp 1597341371
transform 1 0 13524 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1597341371
transform 1 0 14076 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1597341371
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_171
timestamp 1597341371
transform 1 0 16836 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1597341371
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_166
timestamp 1597341371
transform 1 0 16376 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_154
timestamp 1597341371
transform 1 0 15272 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1597341371
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1597341371
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1597341371
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_190
timestamp 1597341371
transform 1 0 18584 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_178
timestamp 1597341371
transform 1 0 17480 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1597341371
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_220
timestamp 1597341371
transform 1 0 21344 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1597341371
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1597341371
transform 1 0 20884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_202
timestamp 1597341371
transform 1 0 19688 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1597341371
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_245
timestamp 1597341371
transform 1 0 23644 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_232
timestamp 1597341371
transform 1 0 22448 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_247
timestamp 1597341371
transform 1 0 23828 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_235
timestamp 1597341371
transform 1 0 22724 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_227
timestamp 1597341371
transform 1 0 21988 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1597341371
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _277_
timestamp 1597341371
transform 1 0 23000 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_47_269
timestamp 1597341371
transform 1 0 25852 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_257
timestamp 1597341371
transform 1 0 24748 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1597341371
transform 1 0 26036 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_259
timestamp 1597341371
transform 1 0 24932 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1597341371
transform 1 0 26956 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_292
timestamp 1597341371
transform 1 0 27968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_288
timestamp 1597341371
transform 1 0 27600 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_276
timestamp 1597341371
transform 1 0 26496 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1597341371
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1597341371
transform -1 0 28336 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1597341371
transform -1 0 28336 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1597341371
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1597341371
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1597341371
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1597341371
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1597341371
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1597341371
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_44
timestamp 1597341371
transform 1 0 5152 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_32
timestamp 1597341371
transform 1 0 4048 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_27
timestamp 1597341371
transform 1 0 3588 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1597341371
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1597341371
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1597341371
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1597341371
transform 1 0 3956 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1597341371
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_63
timestamp 1597341371
transform 1 0 6900 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_56
timestamp 1597341371
transform 1 0 6256 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1597341371
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1597341371
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1597341371
transform 1 0 6808 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1597341371
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_87
timestamp 1597341371
transform 1 0 9108 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_75
timestamp 1597341371
transform 1 0 8004 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1597341371
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1597341371
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1597341371
transform 1 0 9660 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1597341371
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_118
timestamp 1597341371
transform 1 0 11960 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_106
timestamp 1597341371
transform 1 0 10856 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1597341371
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1597341371
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1597341371
transform 1 0 12512 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1597341371
transform 1 0 14812 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1597341371
transform 1 0 13708 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1597341371
transform 1 0 12604 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1597341371
transform 1 0 14076 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1597341371
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_168
timestamp 1597341371
transform 1 0 16560 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_156
timestamp 1597341371
transform 1 0 15456 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1597341371
transform 1 0 16376 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1597341371
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1597341371
transform 1 0 15364 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1597341371
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_187
timestamp 1597341371
transform 1 0 18308 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_180
timestamp 1597341371
transform 1 0 17664 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_190
timestamp 1597341371
transform 1 0 18584 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1597341371
transform 1 0 17480 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1597341371
transform 1 0 18216 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_218
timestamp 1597341371
transform 1 0 21160 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_211
timestamp 1597341371
transform 1 0 20516 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_199
timestamp 1597341371
transform 1 0 19412 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1597341371
transform 1 0 20884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_202
timestamp 1597341371
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1597341371
transform 1 0 21068 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1597341371
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_242
timestamp 1597341371
transform 1 0 23368 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_230
timestamp 1597341371
transform 1 0 22264 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1597341371
transform 1 0 23092 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1597341371
transform 1 0 21988 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1597341371
transform 1 0 23920 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1597341371
transform 1 0 26220 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1597341371
transform 1 0 25116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1597341371
transform 1 0 24012 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_263
timestamp 1597341371
transform 1 0 25300 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_251
timestamp 1597341371
transform 1 0 24196 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_292
timestamp 1597341371
transform 1 0 27968 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_280
timestamp 1597341371
transform 1 0 26864 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_292
timestamp 1597341371
transform 1 0 27968 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_288
timestamp 1597341371
transform 1 0 27600 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_276
timestamp 1597341371
transform 1 0 26496 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1597341371
transform 1 0 26772 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1597341371
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1597341371
transform -1 0 28336 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1597341371
transform -1 0 28336 0 -1 28832
box -38 -48 314 592
<< labels >>
rlabel metal2 s 18510 0 18566 800 6 CSB
port 0 nsew default input
rlabel metal2 s 24858 30864 24914 31664 6 RST
port 1 nsew default input
rlabel metal2 s 9218 0 9274 800 6 SCK
port 2 nsew default input
rlabel metal2 s 18 0 74 800 6 SDI
port 3 nsew default input
rlabel metal3 s 28720 24624 29520 24744 6 mask_rev_in[0]
port 4 nsew default input
rlabel metal3 s 0 27344 800 27464 6 mask_rev_in[1]
port 5 nsew default input
rlabel metal2 s 6366 30864 6422 31664 6 mask_rev_in[2]
port 6 nsew default input
rlabel metal2 s 27710 0 27766 800 6 mask_rev_in[3]
port 7 nsew default input
rlabel metal3 s 28720 11024 29520 11144 6 out
port 8 nsew default tristate
rlabel metal3 s 0 13608 800 13728 6 select
port 9 nsew default input
rlabel metal2 s 15658 30864 15714 31664 6 trap
port 10 nsew default input
rlabel metal5 s 1104 2768 28336 3088 6 VPWR
port 11 nsew default input
rlabel metal5 s 1104 4268 28336 4588 6 VGND
port 12 nsew default input
<< properties >>
string FIXED_BBOX 0 0 29520 31664
<< end >>
